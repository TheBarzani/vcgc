module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 ;
  assign n16 = x3 ^ x0 ;
  assign n17 = x4 ^ x1 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = x5 ^ x2 ;
  assign n20 = n18 & ~n19 ;
  assign n21 = x6 ^ x0 ;
  assign n22 = x7 ^ x1 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = x8 ^ x2 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = ~n20 & ~n25 ;
  assign n27 = x9 ^ x0 ;
  assign n28 = x10 ^ x1 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = x11 ^ x2 ;
  assign n31 = n29 & ~n30 ;
  assign n32 = n26 & ~n31 ;
  assign n33 = x12 ^ x0 ;
  assign n34 = x13 ^ x1 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = x14 ^ x2 ;
  assign n37 = n35 & ~n36 ;
  assign n38 = n32 & ~n37 ;
  assign n39 = x6 ^ x3 ;
  assign n40 = x7 ^ x4 ;
  assign n41 = ~n39 & ~n40 ;
  assign n42 = x8 ^ x5 ;
  assign n43 = n41 & ~n42 ;
  assign n44 = n38 & ~n43 ;
  assign n45 = x9 ^ x3 ;
  assign n46 = x10 ^ x4 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = x11 ^ x5 ;
  assign n49 = n47 & ~n48 ;
  assign n50 = n44 & ~n49 ;
  assign n51 = x12 ^ x3 ;
  assign n52 = x13 ^ x4 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = x14 ^ x5 ;
  assign n55 = n53 & ~n54 ;
  assign n56 = n50 & ~n55 ;
  assign n57 = x9 ^ x6 ;
  assign n58 = x10 ^ x7 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = x11 ^ x8 ;
  assign n61 = n59 & ~n60 ;
  assign n62 = n56 & ~n61 ;
  assign n63 = x12 ^ x6 ;
  assign n64 = x13 ^ x7 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = x14 ^ x8 ;
  assign n67 = n65 & ~n66 ;
  assign n68 = n62 & ~n67 ;
  assign n69 = x12 ^ x9 ;
  assign n70 = x13 ^ x10 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = x14 ^ x11 ;
  assign n73 = n71 & ~n72 ;
  assign n74 = n68 & ~n73 ;
  assign y0 = n74 ;
endmodule
