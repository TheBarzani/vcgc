module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 ;
  output y0 ;
  wire n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 ;
  assign n75 = x2 ^ x0 ;
  assign n76 = x3 ^ x1 ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = x6 ^ x0 ;
  assign n79 = x7 ^ x1 ;
  assign n80 = ~n78 & ~n79 ;
  assign n81 = ~n77 & ~n80 ;
  assign n82 = x20 ^ x0 ;
  assign n83 = x21 ^ x1 ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = n81 & ~n84 ;
  assign n86 = x24 ^ x0 ;
  assign n87 = x25 ^ x1 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = n85 & ~n88 ;
  assign n90 = x4 ^ x2 ;
  assign n91 = x5 ^ x3 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = n89 & ~n92 ;
  assign n94 = x18 ^ x2 ;
  assign n95 = x19 ^ x3 ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = n93 & ~n96 ;
  assign n98 = x22 ^ x2 ;
  assign n99 = x23 ^ x3 ;
  assign n100 = ~n98 & ~n99 ;
  assign n101 = n97 & ~n100 ;
  assign n102 = x10 ^ x4 ;
  assign n103 = x11 ^ x5 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = n101 & ~n104 ;
  assign n106 = x20 ^ x4 ;
  assign n107 = x21 ^ x5 ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = n105 & ~n108 ;
  assign n110 = x28 ^ x4 ;
  assign n111 = x29 ^ x5 ;
  assign n112 = ~n110 & ~n111 ;
  assign n113 = n109 & ~n112 ;
  assign n114 = x8 ^ x6 ;
  assign n115 = x9 ^ x7 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = n113 & ~n116 ;
  assign n118 = x18 ^ x6 ;
  assign n119 = x19 ^ x7 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = n117 & ~n120 ;
  assign n122 = x26 ^ x6 ;
  assign n123 = x27 ^ x7 ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = n121 & ~n124 ;
  assign n126 = x14 ^ x8 ;
  assign n127 = x15 ^ x9 ;
  assign n128 = ~n126 & ~n127 ;
  assign n129 = n125 & ~n128 ;
  assign n130 = x24 ^ x8 ;
  assign n131 = x25 ^ x9 ;
  assign n132 = ~n130 & ~n131 ;
  assign n133 = n129 & ~n132 ;
  assign n134 = x32 ^ x8 ;
  assign n135 = x33 ^ x9 ;
  assign n136 = ~n134 & ~n135 ;
  assign n137 = n133 & ~n136 ;
  assign n138 = x12 ^ x10 ;
  assign n139 = x13 ^ x11 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = n137 & ~n140 ;
  assign n142 = x22 ^ x10 ;
  assign n143 = x23 ^ x11 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = n141 & ~n144 ;
  assign n146 = x30 ^ x10 ;
  assign n147 = x31 ^ x11 ;
  assign n148 = ~n146 & ~n147 ;
  assign n149 = n145 & ~n148 ;
  assign n150 = x16 ^ x12 ;
  assign n151 = x17 ^ x13 ;
  assign n152 = ~n150 & ~n151 ;
  assign n153 = n149 & ~n152 ;
  assign n154 = x28 ^ x12 ;
  assign n155 = x29 ^ x13 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = n153 & ~n156 ;
  assign n158 = x34 ^ x12 ;
  assign n159 = x35 ^ x13 ;
  assign n160 = ~n158 & ~n159 ;
  assign n161 = n157 & ~n160 ;
  assign n162 = x16 ^ x14 ;
  assign n163 = x17 ^ x15 ;
  assign n164 = ~n162 & ~n163 ;
  assign n165 = n161 & ~n164 ;
  assign n166 = x26 ^ x14 ;
  assign n167 = x27 ^ x15 ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = n165 & ~n168 ;
  assign n170 = x34 ^ x14 ;
  assign n171 = x35 ^ x15 ;
  assign n172 = ~n170 & ~n171 ;
  assign n173 = n169 & ~n172 ;
  assign n174 = x30 ^ x16 ;
  assign n175 = x31 ^ x17 ;
  assign n176 = ~n174 & ~n175 ;
  assign n177 = n173 & ~n176 ;
  assign n178 = x32 ^ x16 ;
  assign n179 = x33 ^ x17 ;
  assign n180 = ~n178 & ~n179 ;
  assign n181 = n177 & ~n180 ;
  assign n182 = x38 ^ x18 ;
  assign n183 = x39 ^ x19 ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = n181 & ~n184 ;
  assign n186 = x42 ^ x18 ;
  assign n187 = x43 ^ x19 ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = n185 & ~n188 ;
  assign n190 = x36 ^ x20 ;
  assign n191 = x37 ^ x21 ;
  assign n192 = ~n190 & ~n191 ;
  assign n193 = n189 & ~n192 ;
  assign n194 = x40 ^ x20 ;
  assign n195 = x41 ^ x21 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = n193 & ~n196 ;
  assign n198 = x38 ^ x22 ;
  assign n199 = x39 ^ x23 ;
  assign n200 = ~n198 & ~n199 ;
  assign n201 = n197 & ~n200 ;
  assign n202 = x46 ^ x22 ;
  assign n203 = x47 ^ x23 ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = n201 & ~n204 ;
  assign n206 = x36 ^ x24 ;
  assign n207 = x37 ^ x25 ;
  assign n208 = ~n206 & ~n207 ;
  assign n209 = n205 & ~n208 ;
  assign n210 = x44 ^ x24 ;
  assign n211 = x45 ^ x25 ;
  assign n212 = ~n210 & ~n211 ;
  assign n213 = n209 & ~n212 ;
  assign n214 = x42 ^ x26 ;
  assign n215 = x43 ^ x27 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = n213 & ~n216 ;
  assign n218 = x50 ^ x26 ;
  assign n219 = x51 ^ x27 ;
  assign n220 = ~n218 & ~n219 ;
  assign n221 = n217 & ~n220 ;
  assign n222 = x40 ^ x28 ;
  assign n223 = x41 ^ x29 ;
  assign n224 = ~n222 & ~n223 ;
  assign n225 = n221 & ~n224 ;
  assign n226 = x48 ^ x28 ;
  assign n227 = x49 ^ x29 ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = n225 & ~n228 ;
  assign n230 = x46 ^ x30 ;
  assign n231 = x47 ^ x31 ;
  assign n232 = ~n230 & ~n231 ;
  assign n233 = n229 & ~n232 ;
  assign n234 = x52 ^ x30 ;
  assign n235 = x53 ^ x31 ;
  assign n236 = ~n234 & ~n235 ;
  assign n237 = n233 & ~n236 ;
  assign n238 = x44 ^ x32 ;
  assign n239 = x45 ^ x33 ;
  assign n240 = ~n238 & ~n239 ;
  assign n241 = n237 & ~n240 ;
  assign n242 = x52 ^ x32 ;
  assign n243 = x53 ^ x33 ;
  assign n244 = ~n242 & ~n243 ;
  assign n245 = n241 & ~n244 ;
  assign n246 = x48 ^ x34 ;
  assign n247 = x49 ^ x35 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = n245 & ~n248 ;
  assign n250 = x50 ^ x34 ;
  assign n251 = x51 ^ x35 ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = n249 & ~n252 ;
  assign n254 = x56 ^ x36 ;
  assign n255 = x57 ^ x37 ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = n253 & ~n256 ;
  assign n258 = x60 ^ x36 ;
  assign n259 = x61 ^ x37 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = n257 & ~n260 ;
  assign n262 = x54 ^ x38 ;
  assign n263 = x55 ^ x39 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = n261 & ~n264 ;
  assign n266 = x58 ^ x38 ;
  assign n267 = x59 ^ x39 ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = n265 & ~n268 ;
  assign n270 = x56 ^ x40 ;
  assign n271 = x57 ^ x41 ;
  assign n272 = ~n270 & ~n271 ;
  assign n273 = n269 & ~n272 ;
  assign n274 = x64 ^ x40 ;
  assign n275 = x65 ^ x41 ;
  assign n276 = ~n274 & ~n275 ;
  assign n277 = n273 & ~n276 ;
  assign n278 = x54 ^ x42 ;
  assign n279 = x55 ^ x43 ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = n277 & ~n280 ;
  assign n282 = x62 ^ x42 ;
  assign n283 = x63 ^ x43 ;
  assign n284 = ~n282 & ~n283 ;
  assign n285 = n281 & ~n284 ;
  assign n286 = x60 ^ x44 ;
  assign n287 = x61 ^ x45 ;
  assign n288 = ~n286 & ~n287 ;
  assign n289 = n285 & ~n288 ;
  assign n290 = x68 ^ x44 ;
  assign n291 = x69 ^ x45 ;
  assign n292 = ~n290 & ~n291 ;
  assign n293 = n289 & ~n292 ;
  assign n294 = x58 ^ x46 ;
  assign n295 = x59 ^ x47 ;
  assign n296 = ~n294 & ~n295 ;
  assign n297 = n293 & ~n296 ;
  assign n298 = x66 ^ x46 ;
  assign n299 = x67 ^ x47 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = n297 & ~n300 ;
  assign n302 = x64 ^ x48 ;
  assign n303 = x65 ^ x49 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = n301 & ~n304 ;
  assign n306 = x70 ^ x48 ;
  assign n307 = x71 ^ x49 ;
  assign n308 = ~n306 & ~n307 ;
  assign n309 = n305 & ~n308 ;
  assign n310 = x62 ^ x50 ;
  assign n311 = x63 ^ x51 ;
  assign n312 = ~n310 & ~n311 ;
  assign n313 = n309 & ~n312 ;
  assign n314 = x70 ^ x50 ;
  assign n315 = x71 ^ x51 ;
  assign n316 = ~n314 & ~n315 ;
  assign n317 = n313 & ~n316 ;
  assign n318 = x66 ^ x52 ;
  assign n319 = x67 ^ x53 ;
  assign n320 = ~n318 & ~n319 ;
  assign n321 = n317 & ~n320 ;
  assign n322 = x68 ^ x52 ;
  assign n323 = x69 ^ x53 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = n321 & ~n324 ;
  assign n326 = x72 ^ x54 ;
  assign n327 = x73 ^ x55 ;
  assign n328 = ~n326 & ~n327 ;
  assign n329 = n325 & ~n328 ;
  assign n330 = x72 ^ x56 ;
  assign n331 = x73 ^ x57 ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = n329 & ~n332 ;
  assign n334 = x72 ^ x58 ;
  assign n335 = x73 ^ x59 ;
  assign n336 = ~n334 & ~n335 ;
  assign n337 = n333 & ~n336 ;
  assign n338 = x72 ^ x60 ;
  assign n339 = x73 ^ x61 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n337 & ~n340 ;
  assign n342 = x72 ^ x62 ;
  assign n343 = x73 ^ x63 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = n341 & ~n344 ;
  assign n346 = x72 ^ x64 ;
  assign n347 = x73 ^ x65 ;
  assign n348 = ~n346 & ~n347 ;
  assign n349 = n345 & ~n348 ;
  assign n350 = x72 ^ x66 ;
  assign n351 = x73 ^ x67 ;
  assign n352 = ~n350 & ~n351 ;
  assign n353 = n349 & ~n352 ;
  assign n354 = x72 ^ x68 ;
  assign n355 = x73 ^ x69 ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = n353 & ~n356 ;
  assign n358 = x72 ^ x70 ;
  assign n359 = x73 ^ x71 ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = n357 & ~n360 ;
  assign y0 = n361 ;
endmodule
