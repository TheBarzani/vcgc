module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 ;
  output y0 ;
  wire n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 ;
  assign n142 = x3 ^ x0 ;
  assign n143 = x4 ^ x1 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = x5 ^ x2 ;
  assign n146 = n144 & ~n145 ;
  assign n147 = x9 ^ x0 ;
  assign n148 = x10 ^ x1 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = x11 ^ x2 ;
  assign n151 = n149 & ~n150 ;
  assign n152 = ~n146 & ~n151 ;
  assign n153 = x18 ^ x0 ;
  assign n154 = x19 ^ x1 ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = x20 ^ x2 ;
  assign n157 = n155 & ~n156 ;
  assign n158 = n152 & ~n157 ;
  assign n159 = x24 ^ x0 ;
  assign n160 = x25 ^ x1 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = x26 ^ x2 ;
  assign n163 = n161 & ~n162 ;
  assign n164 = n158 & ~n163 ;
  assign n165 = x36 ^ x0 ;
  assign n166 = x37 ^ x1 ;
  assign n167 = ~n165 & ~n166 ;
  assign n168 = x38 ^ x2 ;
  assign n169 = n167 & ~n168 ;
  assign n170 = n164 & ~n169 ;
  assign n171 = x42 ^ x0 ;
  assign n172 = x43 ^ x1 ;
  assign n173 = ~n171 & ~n172 ;
  assign n174 = x44 ^ x2 ;
  assign n175 = n173 & ~n174 ;
  assign n176 = n170 & ~n175 ;
  assign n177 = x51 ^ x0 ;
  assign n178 = x52 ^ x1 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = x53 ^ x2 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n176 & ~n181 ;
  assign n183 = x57 ^ x0 ;
  assign n184 = x58 ^ x1 ;
  assign n185 = ~n183 & ~n184 ;
  assign n186 = x59 ^ x2 ;
  assign n187 = n185 & ~n186 ;
  assign n188 = n182 & ~n187 ;
  assign n189 = x72 ^ x0 ;
  assign n190 = x73 ^ x1 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = x74 ^ x2 ;
  assign n193 = n191 & ~n192 ;
  assign n194 = n188 & ~n193 ;
  assign n195 = x78 ^ x0 ;
  assign n196 = x79 ^ x1 ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = x80 ^ x2 ;
  assign n199 = n197 & ~n198 ;
  assign n200 = n194 & ~n199 ;
  assign n201 = x87 ^ x0 ;
  assign n202 = x88 ^ x1 ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = x89 ^ x2 ;
  assign n205 = n203 & ~n204 ;
  assign n206 = n200 & ~n205 ;
  assign n207 = x93 ^ x0 ;
  assign n208 = x94 ^ x1 ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = x95 ^ x2 ;
  assign n211 = n209 & ~n210 ;
  assign n212 = n206 & ~n211 ;
  assign n213 = x105 ^ x0 ;
  assign n214 = x106 ^ x1 ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = x107 ^ x2 ;
  assign n217 = n215 & ~n216 ;
  assign n218 = n212 & ~n217 ;
  assign n219 = x111 ^ x0 ;
  assign n220 = x112 ^ x1 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = x113 ^ x2 ;
  assign n223 = n221 & ~n222 ;
  assign n224 = n218 & ~n223 ;
  assign n225 = x120 ^ x0 ;
  assign n226 = x121 ^ x1 ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = x122 ^ x2 ;
  assign n229 = n227 & ~n228 ;
  assign n230 = n224 & ~n229 ;
  assign n231 = x126 ^ x0 ;
  assign n232 = x127 ^ x1 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = x128 ^ x2 ;
  assign n235 = n233 & ~n234 ;
  assign n236 = n230 & ~n235 ;
  assign n237 = x6 ^ x3 ;
  assign n238 = x7 ^ x4 ;
  assign n239 = ~n237 & ~n238 ;
  assign n240 = x8 ^ x5 ;
  assign n241 = n239 & ~n240 ;
  assign n242 = n236 & ~n241 ;
  assign n243 = x15 ^ x3 ;
  assign n244 = x16 ^ x4 ;
  assign n245 = ~n243 & ~n244 ;
  assign n246 = x17 ^ x5 ;
  assign n247 = n245 & ~n246 ;
  assign n248 = n242 & ~n247 ;
  assign n249 = x21 ^ x3 ;
  assign n250 = x22 ^ x4 ;
  assign n251 = ~n249 & ~n250 ;
  assign n252 = x23 ^ x5 ;
  assign n253 = n251 & ~n252 ;
  assign n254 = n248 & ~n253 ;
  assign n255 = x33 ^ x3 ;
  assign n256 = x34 ^ x4 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = x35 ^ x5 ;
  assign n259 = n257 & ~n258 ;
  assign n260 = n254 & ~n259 ;
  assign n261 = x39 ^ x3 ;
  assign n262 = x40 ^ x4 ;
  assign n263 = ~n261 & ~n262 ;
  assign n264 = x41 ^ x5 ;
  assign n265 = n263 & ~n264 ;
  assign n266 = n260 & ~n265 ;
  assign n267 = x48 ^ x3 ;
  assign n268 = x49 ^ x4 ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = x50 ^ x5 ;
  assign n271 = n269 & ~n270 ;
  assign n272 = n266 & ~n271 ;
  assign n273 = x54 ^ x3 ;
  assign n274 = x55 ^ x4 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = x56 ^ x5 ;
  assign n277 = n275 & ~n276 ;
  assign n278 = n272 & ~n277 ;
  assign n279 = x69 ^ x3 ;
  assign n280 = x70 ^ x4 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = x71 ^ x5 ;
  assign n283 = n281 & ~n282 ;
  assign n284 = n278 & ~n283 ;
  assign n285 = x75 ^ x3 ;
  assign n286 = x76 ^ x4 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = x77 ^ x5 ;
  assign n289 = n287 & ~n288 ;
  assign n290 = n284 & ~n289 ;
  assign n291 = x84 ^ x3 ;
  assign n292 = x85 ^ x4 ;
  assign n293 = ~n291 & ~n292 ;
  assign n294 = x86 ^ x5 ;
  assign n295 = n293 & ~n294 ;
  assign n296 = n290 & ~n295 ;
  assign n297 = x90 ^ x3 ;
  assign n298 = x91 ^ x4 ;
  assign n299 = ~n297 & ~n298 ;
  assign n300 = x92 ^ x5 ;
  assign n301 = n299 & ~n300 ;
  assign n302 = n296 & ~n301 ;
  assign n303 = x102 ^ x3 ;
  assign n304 = x103 ^ x4 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = x104 ^ x5 ;
  assign n307 = n305 & ~n306 ;
  assign n308 = n302 & ~n307 ;
  assign n309 = x108 ^ x3 ;
  assign n310 = x109 ^ x4 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = x110 ^ x5 ;
  assign n313 = n311 & ~n312 ;
  assign n314 = n308 & ~n313 ;
  assign n315 = x117 ^ x3 ;
  assign n316 = x118 ^ x4 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = x119 ^ x5 ;
  assign n319 = n317 & ~n318 ;
  assign n320 = n314 & ~n319 ;
  assign n321 = x123 ^ x3 ;
  assign n322 = x124 ^ x4 ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = x125 ^ x5 ;
  assign n325 = n323 & ~n324 ;
  assign n326 = n320 & ~n325 ;
  assign n327 = x12 ^ x6 ;
  assign n328 = x13 ^ x7 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = x14 ^ x8 ;
  assign n331 = n329 & ~n330 ;
  assign n332 = n326 & ~n331 ;
  assign n333 = x18 ^ x6 ;
  assign n334 = x19 ^ x7 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = x20 ^ x8 ;
  assign n337 = n335 & ~n336 ;
  assign n338 = n332 & ~n337 ;
  assign n339 = x27 ^ x6 ;
  assign n340 = x28 ^ x7 ;
  assign n341 = ~n339 & ~n340 ;
  assign n342 = x29 ^ x8 ;
  assign n343 = n341 & ~n342 ;
  assign n344 = n338 & ~n343 ;
  assign n345 = x36 ^ x6 ;
  assign n346 = x37 ^ x7 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = x38 ^ x8 ;
  assign n349 = n347 & ~n348 ;
  assign n350 = n344 & ~n349 ;
  assign n351 = x45 ^ x6 ;
  assign n352 = x46 ^ x7 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = x47 ^ x8 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = n350 & ~n355 ;
  assign n357 = x51 ^ x6 ;
  assign n358 = x52 ^ x7 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = x53 ^ x8 ;
  assign n361 = n359 & ~n360 ;
  assign n362 = n356 & ~n361 ;
  assign n363 = x60 ^ x6 ;
  assign n364 = x61 ^ x7 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = x62 ^ x8 ;
  assign n367 = n365 & ~n366 ;
  assign n368 = n362 & ~n367 ;
  assign n369 = x72 ^ x6 ;
  assign n370 = x73 ^ x7 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = x74 ^ x8 ;
  assign n373 = n371 & ~n372 ;
  assign n374 = n368 & ~n373 ;
  assign n375 = x81 ^ x6 ;
  assign n376 = x82 ^ x7 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = x83 ^ x8 ;
  assign n379 = n377 & ~n378 ;
  assign n380 = n374 & ~n379 ;
  assign n381 = x87 ^ x6 ;
  assign n382 = x88 ^ x7 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = x89 ^ x8 ;
  assign n385 = n383 & ~n384 ;
  assign n386 = n380 & ~n385 ;
  assign n387 = x96 ^ x6 ;
  assign n388 = x97 ^ x7 ;
  assign n389 = ~n387 & ~n388 ;
  assign n390 = x98 ^ x8 ;
  assign n391 = n389 & ~n390 ;
  assign n392 = n386 & ~n391 ;
  assign n393 = x105 ^ x6 ;
  assign n394 = x106 ^ x7 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = x107 ^ x8 ;
  assign n397 = n395 & ~n396 ;
  assign n398 = n392 & ~n397 ;
  assign n399 = x114 ^ x6 ;
  assign n400 = x115 ^ x7 ;
  assign n401 = ~n399 & ~n400 ;
  assign n402 = x116 ^ x8 ;
  assign n403 = n401 & ~n402 ;
  assign n404 = n398 & ~n403 ;
  assign n405 = x120 ^ x6 ;
  assign n406 = x121 ^ x7 ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = x122 ^ x8 ;
  assign n409 = n407 & ~n408 ;
  assign n410 = n404 & ~n409 ;
  assign n411 = x129 ^ x6 ;
  assign n412 = x130 ^ x7 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = x131 ^ x8 ;
  assign n415 = n413 & ~n414 ;
  assign n416 = n410 & ~n415 ;
  assign n417 = x12 ^ x9 ;
  assign n418 = x13 ^ x10 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = x14 ^ x11 ;
  assign n421 = n419 & ~n420 ;
  assign n422 = n416 & ~n421 ;
  assign n423 = x15 ^ x9 ;
  assign n424 = x16 ^ x10 ;
  assign n425 = ~n423 & ~n424 ;
  assign n426 = x17 ^ x11 ;
  assign n427 = n425 & ~n426 ;
  assign n428 = n422 & ~n427 ;
  assign n429 = x27 ^ x9 ;
  assign n430 = x28 ^ x10 ;
  assign n431 = ~n429 & ~n430 ;
  assign n432 = x29 ^ x11 ;
  assign n433 = n431 & ~n432 ;
  assign n434 = n428 & ~n433 ;
  assign n435 = x33 ^ x9 ;
  assign n436 = x34 ^ x10 ;
  assign n437 = ~n435 & ~n436 ;
  assign n438 = x35 ^ x11 ;
  assign n439 = n437 & ~n438 ;
  assign n440 = n434 & ~n439 ;
  assign n441 = x45 ^ x9 ;
  assign n442 = x46 ^ x10 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = x47 ^ x11 ;
  assign n445 = n443 & ~n444 ;
  assign n446 = n440 & ~n445 ;
  assign n447 = x48 ^ x9 ;
  assign n448 = x49 ^ x10 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = x50 ^ x11 ;
  assign n451 = n449 & ~n450 ;
  assign n452 = n446 & ~n451 ;
  assign n453 = x60 ^ x9 ;
  assign n454 = x61 ^ x10 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = x62 ^ x11 ;
  assign n457 = n455 & ~n456 ;
  assign n458 = n452 & ~n457 ;
  assign n459 = x69 ^ x9 ;
  assign n460 = x70 ^ x10 ;
  assign n461 = ~n459 & ~n460 ;
  assign n462 = x71 ^ x11 ;
  assign n463 = n461 & ~n462 ;
  assign n464 = n458 & ~n463 ;
  assign n465 = x81 ^ x9 ;
  assign n466 = x82 ^ x10 ;
  assign n467 = ~n465 & ~n466 ;
  assign n468 = x83 ^ x11 ;
  assign n469 = n467 & ~n468 ;
  assign n470 = n464 & ~n469 ;
  assign n471 = x84 ^ x9 ;
  assign n472 = x85 ^ x10 ;
  assign n473 = ~n471 & ~n472 ;
  assign n474 = x86 ^ x11 ;
  assign n475 = n473 & ~n474 ;
  assign n476 = n470 & ~n475 ;
  assign n477 = x96 ^ x9 ;
  assign n478 = x97 ^ x10 ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = x98 ^ x11 ;
  assign n481 = n479 & ~n480 ;
  assign n482 = n476 & ~n481 ;
  assign n483 = x102 ^ x9 ;
  assign n484 = x103 ^ x10 ;
  assign n485 = ~n483 & ~n484 ;
  assign n486 = x104 ^ x11 ;
  assign n487 = n485 & ~n486 ;
  assign n488 = n482 & ~n487 ;
  assign n489 = x114 ^ x9 ;
  assign n490 = x115 ^ x10 ;
  assign n491 = ~n489 & ~n490 ;
  assign n492 = x116 ^ x11 ;
  assign n493 = n491 & ~n492 ;
  assign n494 = n488 & ~n493 ;
  assign n495 = x117 ^ x9 ;
  assign n496 = x118 ^ x10 ;
  assign n497 = ~n495 & ~n496 ;
  assign n498 = x119 ^ x11 ;
  assign n499 = n497 & ~n498 ;
  assign n500 = n494 & ~n499 ;
  assign n501 = x129 ^ x9 ;
  assign n502 = x130 ^ x10 ;
  assign n503 = ~n501 & ~n502 ;
  assign n504 = x131 ^ x11 ;
  assign n505 = n503 & ~n504 ;
  assign n506 = n500 & ~n505 ;
  assign n507 = x21 ^ x12 ;
  assign n508 = x22 ^ x13 ;
  assign n509 = ~n507 & ~n508 ;
  assign n510 = x23 ^ x14 ;
  assign n511 = n509 & ~n510 ;
  assign n512 = n506 & ~n511 ;
  assign n513 = x24 ^ x12 ;
  assign n514 = x25 ^ x13 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = x26 ^ x14 ;
  assign n517 = n515 & ~n516 ;
  assign n518 = n512 & ~n517 ;
  assign n519 = x39 ^ x12 ;
  assign n520 = x40 ^ x13 ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = x41 ^ x14 ;
  assign n523 = n521 & ~n522 ;
  assign n524 = n518 & ~n523 ;
  assign n525 = x42 ^ x12 ;
  assign n526 = x43 ^ x13 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = x44 ^ x14 ;
  assign n529 = n527 & ~n528 ;
  assign n530 = n524 & ~n529 ;
  assign n531 = x54 ^ x12 ;
  assign n532 = x55 ^ x13 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = x56 ^ x14 ;
  assign n535 = n533 & ~n534 ;
  assign n536 = n530 & ~n535 ;
  assign n537 = x57 ^ x12 ;
  assign n538 = x58 ^ x13 ;
  assign n539 = ~n537 & ~n538 ;
  assign n540 = x59 ^ x14 ;
  assign n541 = n539 & ~n540 ;
  assign n542 = n536 & ~n541 ;
  assign n543 = x75 ^ x12 ;
  assign n544 = x76 ^ x13 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = x77 ^ x14 ;
  assign n547 = n545 & ~n546 ;
  assign n548 = n542 & ~n547 ;
  assign n549 = x78 ^ x12 ;
  assign n550 = x79 ^ x13 ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = x80 ^ x14 ;
  assign n553 = n551 & ~n552 ;
  assign n554 = n548 & ~n553 ;
  assign n555 = x90 ^ x12 ;
  assign n556 = x91 ^ x13 ;
  assign n557 = ~n555 & ~n556 ;
  assign n558 = x92 ^ x14 ;
  assign n559 = n557 & ~n558 ;
  assign n560 = n554 & ~n559 ;
  assign n561 = x93 ^ x12 ;
  assign n562 = x94 ^ x13 ;
  assign n563 = ~n561 & ~n562 ;
  assign n564 = x95 ^ x14 ;
  assign n565 = n563 & ~n564 ;
  assign n566 = n560 & ~n565 ;
  assign n567 = x108 ^ x12 ;
  assign n568 = x109 ^ x13 ;
  assign n569 = ~n567 & ~n568 ;
  assign n570 = x110 ^ x14 ;
  assign n571 = n569 & ~n570 ;
  assign n572 = n566 & ~n571 ;
  assign n573 = x111 ^ x12 ;
  assign n574 = x112 ^ x13 ;
  assign n575 = ~n573 & ~n574 ;
  assign n576 = x113 ^ x14 ;
  assign n577 = n575 & ~n576 ;
  assign n578 = n572 & ~n577 ;
  assign n579 = x123 ^ x12 ;
  assign n580 = x124 ^ x13 ;
  assign n581 = ~n579 & ~n580 ;
  assign n582 = x125 ^ x14 ;
  assign n583 = n581 & ~n582 ;
  assign n584 = n578 & ~n583 ;
  assign n585 = x126 ^ x12 ;
  assign n586 = x127 ^ x13 ;
  assign n587 = ~n585 & ~n586 ;
  assign n588 = x128 ^ x14 ;
  assign n589 = n587 & ~n588 ;
  assign n590 = n584 & ~n589 ;
  assign n591 = x30 ^ x15 ;
  assign n592 = x31 ^ x16 ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = x32 ^ x17 ;
  assign n595 = n593 & ~n594 ;
  assign n596 = n590 & ~n595 ;
  assign n597 = x36 ^ x15 ;
  assign n598 = x37 ^ x16 ;
  assign n599 = ~n597 & ~n598 ;
  assign n600 = x38 ^ x17 ;
  assign n601 = n599 & ~n600 ;
  assign n602 = n596 & ~n601 ;
  assign n603 = x42 ^ x15 ;
  assign n604 = x43 ^ x16 ;
  assign n605 = ~n603 & ~n604 ;
  assign n606 = x44 ^ x17 ;
  assign n607 = n605 & ~n606 ;
  assign n608 = n602 & ~n607 ;
  assign n609 = x63 ^ x15 ;
  assign n610 = x64 ^ x16 ;
  assign n611 = ~n609 & ~n610 ;
  assign n612 = x65 ^ x17 ;
  assign n613 = n611 & ~n612 ;
  assign n614 = n608 & ~n613 ;
  assign n615 = x72 ^ x15 ;
  assign n616 = x73 ^ x16 ;
  assign n617 = ~n615 & ~n616 ;
  assign n618 = x74 ^ x17 ;
  assign n619 = n617 & ~n618 ;
  assign n620 = n614 & ~n619 ;
  assign n621 = x78 ^ x15 ;
  assign n622 = x79 ^ x16 ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = x80 ^ x17 ;
  assign n625 = n623 & ~n624 ;
  assign n626 = n620 & ~n625 ;
  assign n627 = x99 ^ x15 ;
  assign n628 = x100 ^ x16 ;
  assign n629 = ~n627 & ~n628 ;
  assign n630 = x101 ^ x17 ;
  assign n631 = n629 & ~n630 ;
  assign n632 = n626 & ~n631 ;
  assign n633 = x105 ^ x15 ;
  assign n634 = x106 ^ x16 ;
  assign n635 = ~n633 & ~n634 ;
  assign n636 = x107 ^ x17 ;
  assign n637 = n635 & ~n636 ;
  assign n638 = n632 & ~n637 ;
  assign n639 = x111 ^ x15 ;
  assign n640 = x112 ^ x16 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = x113 ^ x17 ;
  assign n643 = n641 & ~n642 ;
  assign n644 = n638 & ~n643 ;
  assign n645 = x132 ^ x15 ;
  assign n646 = x133 ^ x16 ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = x134 ^ x17 ;
  assign n649 = n647 & ~n648 ;
  assign n650 = n644 & ~n649 ;
  assign n651 = x30 ^ x18 ;
  assign n652 = x31 ^ x19 ;
  assign n653 = ~n651 & ~n652 ;
  assign n654 = x32 ^ x20 ;
  assign n655 = n653 & ~n654 ;
  assign n656 = n650 & ~n655 ;
  assign n657 = x33 ^ x18 ;
  assign n658 = x34 ^ x19 ;
  assign n659 = ~n657 & ~n658 ;
  assign n660 = x35 ^ x20 ;
  assign n661 = n659 & ~n660 ;
  assign n662 = n656 & ~n661 ;
  assign n663 = x39 ^ x18 ;
  assign n664 = x40 ^ x19 ;
  assign n665 = ~n663 & ~n664 ;
  assign n666 = x41 ^ x20 ;
  assign n667 = n665 & ~n666 ;
  assign n668 = n662 & ~n667 ;
  assign n669 = x63 ^ x18 ;
  assign n670 = x64 ^ x19 ;
  assign n671 = ~n669 & ~n670 ;
  assign n672 = x65 ^ x20 ;
  assign n673 = n671 & ~n672 ;
  assign n674 = n668 & ~n673 ;
  assign n675 = x69 ^ x18 ;
  assign n676 = x70 ^ x19 ;
  assign n677 = ~n675 & ~n676 ;
  assign n678 = x71 ^ x20 ;
  assign n679 = n677 & ~n678 ;
  assign n680 = n674 & ~n679 ;
  assign n681 = x75 ^ x18 ;
  assign n682 = x76 ^ x19 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = x77 ^ x20 ;
  assign n685 = n683 & ~n684 ;
  assign n686 = n680 & ~n685 ;
  assign n687 = x99 ^ x18 ;
  assign n688 = x100 ^ x19 ;
  assign n689 = ~n687 & ~n688 ;
  assign n690 = x101 ^ x20 ;
  assign n691 = n689 & ~n690 ;
  assign n692 = n686 & ~n691 ;
  assign n693 = x102 ^ x18 ;
  assign n694 = x103 ^ x19 ;
  assign n695 = ~n693 & ~n694 ;
  assign n696 = x104 ^ x20 ;
  assign n697 = n695 & ~n696 ;
  assign n698 = n692 & ~n697 ;
  assign n699 = x108 ^ x18 ;
  assign n700 = x109 ^ x19 ;
  assign n701 = ~n699 & ~n700 ;
  assign n702 = x110 ^ x20 ;
  assign n703 = n701 & ~n702 ;
  assign n704 = n698 & ~n703 ;
  assign n705 = x132 ^ x18 ;
  assign n706 = x133 ^ x19 ;
  assign n707 = ~n705 & ~n706 ;
  assign n708 = x134 ^ x20 ;
  assign n709 = n707 & ~n708 ;
  assign n710 = n704 & ~n709 ;
  assign n711 = x30 ^ x21 ;
  assign n712 = x31 ^ x22 ;
  assign n713 = ~n711 & ~n712 ;
  assign n714 = x32 ^ x23 ;
  assign n715 = n713 & ~n714 ;
  assign n716 = n710 & ~n715 ;
  assign n717 = x36 ^ x21 ;
  assign n718 = x37 ^ x22 ;
  assign n719 = ~n717 & ~n718 ;
  assign n720 = x38 ^ x23 ;
  assign n721 = n719 & ~n720 ;
  assign n722 = n716 & ~n721 ;
  assign n723 = x45 ^ x21 ;
  assign n724 = x46 ^ x22 ;
  assign n725 = ~n723 & ~n724 ;
  assign n726 = x47 ^ x23 ;
  assign n727 = n725 & ~n726 ;
  assign n728 = n722 & ~n727 ;
  assign n729 = x63 ^ x21 ;
  assign n730 = x64 ^ x22 ;
  assign n731 = ~n729 & ~n730 ;
  assign n732 = x65 ^ x23 ;
  assign n733 = n731 & ~n732 ;
  assign n734 = n728 & ~n733 ;
  assign n735 = x72 ^ x21 ;
  assign n736 = x73 ^ x22 ;
  assign n737 = ~n735 & ~n736 ;
  assign n738 = x74 ^ x23 ;
  assign n739 = n737 & ~n738 ;
  assign n740 = n734 & ~n739 ;
  assign n741 = x81 ^ x21 ;
  assign n742 = x82 ^ x22 ;
  assign n743 = ~n741 & ~n742 ;
  assign n744 = x83 ^ x23 ;
  assign n745 = n743 & ~n744 ;
  assign n746 = n740 & ~n745 ;
  assign n747 = x99 ^ x21 ;
  assign n748 = x100 ^ x22 ;
  assign n749 = ~n747 & ~n748 ;
  assign n750 = x101 ^ x23 ;
  assign n751 = n749 & ~n750 ;
  assign n752 = n746 & ~n751 ;
  assign n753 = x105 ^ x21 ;
  assign n754 = x106 ^ x22 ;
  assign n755 = ~n753 & ~n754 ;
  assign n756 = x107 ^ x23 ;
  assign n757 = n755 & ~n756 ;
  assign n758 = n752 & ~n757 ;
  assign n759 = x114 ^ x21 ;
  assign n760 = x115 ^ x22 ;
  assign n761 = ~n759 & ~n760 ;
  assign n762 = x116 ^ x23 ;
  assign n763 = n761 & ~n762 ;
  assign n764 = n758 & ~n763 ;
  assign n765 = x132 ^ x21 ;
  assign n766 = x133 ^ x22 ;
  assign n767 = ~n765 & ~n766 ;
  assign n768 = x134 ^ x23 ;
  assign n769 = n767 & ~n768 ;
  assign n770 = n764 & ~n769 ;
  assign n771 = x30 ^ x24 ;
  assign n772 = x31 ^ x25 ;
  assign n773 = ~n771 & ~n772 ;
  assign n774 = x32 ^ x26 ;
  assign n775 = n773 & ~n774 ;
  assign n776 = n770 & ~n775 ;
  assign n777 = x33 ^ x24 ;
  assign n778 = x34 ^ x25 ;
  assign n779 = ~n777 & ~n778 ;
  assign n780 = x35 ^ x26 ;
  assign n781 = n779 & ~n780 ;
  assign n782 = n776 & ~n781 ;
  assign n783 = x45 ^ x24 ;
  assign n784 = x46 ^ x25 ;
  assign n785 = ~n783 & ~n784 ;
  assign n786 = x47 ^ x26 ;
  assign n787 = n785 & ~n786 ;
  assign n788 = n782 & ~n787 ;
  assign n789 = x63 ^ x24 ;
  assign n790 = x64 ^ x25 ;
  assign n791 = ~n789 & ~n790 ;
  assign n792 = x65 ^ x26 ;
  assign n793 = n791 & ~n792 ;
  assign n794 = n788 & ~n793 ;
  assign n795 = x69 ^ x24 ;
  assign n796 = x70 ^ x25 ;
  assign n797 = ~n795 & ~n796 ;
  assign n798 = x71 ^ x26 ;
  assign n799 = n797 & ~n798 ;
  assign n800 = n794 & ~n799 ;
  assign n801 = x81 ^ x24 ;
  assign n802 = x82 ^ x25 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = x83 ^ x26 ;
  assign n805 = n803 & ~n804 ;
  assign n806 = n800 & ~n805 ;
  assign n807 = x99 ^ x24 ;
  assign n808 = x100 ^ x25 ;
  assign n809 = ~n807 & ~n808 ;
  assign n810 = x101 ^ x26 ;
  assign n811 = n809 & ~n810 ;
  assign n812 = n806 & ~n811 ;
  assign n813 = x102 ^ x24 ;
  assign n814 = x103 ^ x25 ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = x104 ^ x26 ;
  assign n817 = n815 & ~n816 ;
  assign n818 = n812 & ~n817 ;
  assign n819 = x114 ^ x24 ;
  assign n820 = x115 ^ x25 ;
  assign n821 = ~n819 & ~n820 ;
  assign n822 = x116 ^ x26 ;
  assign n823 = n821 & ~n822 ;
  assign n824 = n818 & ~n823 ;
  assign n825 = x132 ^ x24 ;
  assign n826 = x133 ^ x25 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = x134 ^ x26 ;
  assign n829 = n827 & ~n828 ;
  assign n830 = n824 & ~n829 ;
  assign n831 = x30 ^ x27 ;
  assign n832 = x31 ^ x28 ;
  assign n833 = ~n831 & ~n832 ;
  assign n834 = x32 ^ x29 ;
  assign n835 = n833 & ~n834 ;
  assign n836 = n830 & ~n835 ;
  assign n837 = x39 ^ x27 ;
  assign n838 = x40 ^ x28 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = x41 ^ x29 ;
  assign n841 = n839 & ~n840 ;
  assign n842 = n836 & ~n841 ;
  assign n843 = x42 ^ x27 ;
  assign n844 = x43 ^ x28 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = x44 ^ x29 ;
  assign n847 = n845 & ~n846 ;
  assign n848 = n842 & ~n847 ;
  assign n849 = x63 ^ x27 ;
  assign n850 = x64 ^ x28 ;
  assign n851 = ~n849 & ~n850 ;
  assign n852 = x65 ^ x29 ;
  assign n853 = n851 & ~n852 ;
  assign n854 = n848 & ~n853 ;
  assign n855 = x75 ^ x27 ;
  assign n856 = x76 ^ x28 ;
  assign n857 = ~n855 & ~n856 ;
  assign n858 = x77 ^ x29 ;
  assign n859 = n857 & ~n858 ;
  assign n860 = n854 & ~n859 ;
  assign n861 = x78 ^ x27 ;
  assign n862 = x79 ^ x28 ;
  assign n863 = ~n861 & ~n862 ;
  assign n864 = x80 ^ x29 ;
  assign n865 = n863 & ~n864 ;
  assign n866 = n860 & ~n865 ;
  assign n867 = x99 ^ x27 ;
  assign n868 = x100 ^ x28 ;
  assign n869 = ~n867 & ~n868 ;
  assign n870 = x101 ^ x29 ;
  assign n871 = n869 & ~n870 ;
  assign n872 = n866 & ~n871 ;
  assign n873 = x108 ^ x27 ;
  assign n874 = x109 ^ x28 ;
  assign n875 = ~n873 & ~n874 ;
  assign n876 = x110 ^ x29 ;
  assign n877 = n875 & ~n876 ;
  assign n878 = n872 & ~n877 ;
  assign n879 = x111 ^ x27 ;
  assign n880 = x112 ^ x28 ;
  assign n881 = ~n879 & ~n880 ;
  assign n882 = x113 ^ x29 ;
  assign n883 = n881 & ~n882 ;
  assign n884 = n878 & ~n883 ;
  assign n885 = x132 ^ x27 ;
  assign n886 = x133 ^ x28 ;
  assign n887 = ~n885 & ~n886 ;
  assign n888 = x134 ^ x29 ;
  assign n889 = n887 & ~n888 ;
  assign n890 = n884 & ~n889 ;
  assign n891 = x48 ^ x30 ;
  assign n892 = x49 ^ x31 ;
  assign n893 = ~n891 & ~n892 ;
  assign n894 = x50 ^ x32 ;
  assign n895 = n893 & ~n894 ;
  assign n896 = n890 & ~n895 ;
  assign n897 = x51 ^ x30 ;
  assign n898 = x52 ^ x31 ;
  assign n899 = ~n897 & ~n898 ;
  assign n900 = x53 ^ x32 ;
  assign n901 = n899 & ~n900 ;
  assign n902 = n896 & ~n901 ;
  assign n903 = x54 ^ x30 ;
  assign n904 = x55 ^ x31 ;
  assign n905 = ~n903 & ~n904 ;
  assign n906 = x56 ^ x32 ;
  assign n907 = n905 & ~n906 ;
  assign n908 = n902 & ~n907 ;
  assign n909 = x57 ^ x30 ;
  assign n910 = x58 ^ x31 ;
  assign n911 = ~n909 & ~n910 ;
  assign n912 = x59 ^ x32 ;
  assign n913 = n911 & ~n912 ;
  assign n914 = n908 & ~n913 ;
  assign n915 = x60 ^ x30 ;
  assign n916 = x61 ^ x31 ;
  assign n917 = ~n915 & ~n916 ;
  assign n918 = x62 ^ x32 ;
  assign n919 = n917 & ~n918 ;
  assign n920 = n914 & ~n919 ;
  assign n921 = x84 ^ x30 ;
  assign n922 = x85 ^ x31 ;
  assign n923 = ~n921 & ~n922 ;
  assign n924 = x86 ^ x32 ;
  assign n925 = n923 & ~n924 ;
  assign n926 = n920 & ~n925 ;
  assign n927 = x87 ^ x30 ;
  assign n928 = x88 ^ x31 ;
  assign n929 = ~n927 & ~n928 ;
  assign n930 = x89 ^ x32 ;
  assign n931 = n929 & ~n930 ;
  assign n932 = n926 & ~n931 ;
  assign n933 = x90 ^ x30 ;
  assign n934 = x91 ^ x31 ;
  assign n935 = ~n933 & ~n934 ;
  assign n936 = x92 ^ x32 ;
  assign n937 = n935 & ~n936 ;
  assign n938 = n932 & ~n937 ;
  assign n939 = x93 ^ x30 ;
  assign n940 = x94 ^ x31 ;
  assign n941 = ~n939 & ~n940 ;
  assign n942 = x95 ^ x32 ;
  assign n943 = n941 & ~n942 ;
  assign n944 = n938 & ~n943 ;
  assign n945 = x96 ^ x30 ;
  assign n946 = x97 ^ x31 ;
  assign n947 = ~n945 & ~n946 ;
  assign n948 = x98 ^ x32 ;
  assign n949 = n947 & ~n948 ;
  assign n950 = n944 & ~n949 ;
  assign n951 = x117 ^ x30 ;
  assign n952 = x118 ^ x31 ;
  assign n953 = ~n951 & ~n952 ;
  assign n954 = x119 ^ x32 ;
  assign n955 = n953 & ~n954 ;
  assign n956 = n950 & ~n955 ;
  assign n957 = x120 ^ x30 ;
  assign n958 = x121 ^ x31 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = x122 ^ x32 ;
  assign n961 = n959 & ~n960 ;
  assign n962 = n956 & ~n961 ;
  assign n963 = x123 ^ x30 ;
  assign n964 = x124 ^ x31 ;
  assign n965 = ~n963 & ~n964 ;
  assign n966 = x125 ^ x32 ;
  assign n967 = n965 & ~n966 ;
  assign n968 = n962 & ~n967 ;
  assign n969 = x126 ^ x30 ;
  assign n970 = x127 ^ x31 ;
  assign n971 = ~n969 & ~n970 ;
  assign n972 = x128 ^ x32 ;
  assign n973 = n971 & ~n972 ;
  assign n974 = n968 & ~n973 ;
  assign n975 = x129 ^ x30 ;
  assign n976 = x130 ^ x31 ;
  assign n977 = ~n975 & ~n976 ;
  assign n978 = x131 ^ x32 ;
  assign n979 = n977 & ~n978 ;
  assign n980 = n974 & ~n979 ;
  assign n981 = x66 ^ x33 ;
  assign n982 = x67 ^ x34 ;
  assign n983 = ~n981 & ~n982 ;
  assign n984 = x68 ^ x35 ;
  assign n985 = n983 & ~n984 ;
  assign n986 = n980 & ~n985 ;
  assign n987 = x72 ^ x33 ;
  assign n988 = x73 ^ x34 ;
  assign n989 = ~n987 & ~n988 ;
  assign n990 = x74 ^ x35 ;
  assign n991 = n989 & ~n990 ;
  assign n992 = n986 & ~n991 ;
  assign n993 = x78 ^ x33 ;
  assign n994 = x79 ^ x34 ;
  assign n995 = ~n993 & ~n994 ;
  assign n996 = x80 ^ x35 ;
  assign n997 = n995 & ~n996 ;
  assign n998 = n992 & ~n997 ;
  assign n999 = x87 ^ x33 ;
  assign n1000 = x88 ^ x34 ;
  assign n1001 = ~n999 & ~n1000 ;
  assign n1002 = x89 ^ x35 ;
  assign n1003 = n1001 & ~n1002 ;
  assign n1004 = n998 & ~n1003 ;
  assign n1005 = x93 ^ x33 ;
  assign n1006 = x94 ^ x34 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = x95 ^ x35 ;
  assign n1009 = n1007 & ~n1008 ;
  assign n1010 = n1004 & ~n1009 ;
  assign n1011 = x135 ^ x33 ;
  assign n1012 = x136 ^ x34 ;
  assign n1013 = ~n1011 & ~n1012 ;
  assign n1014 = x137 ^ x35 ;
  assign n1015 = n1013 & ~n1014 ;
  assign n1016 = n1010 & ~n1015 ;
  assign n1017 = x66 ^ x36 ;
  assign n1018 = x67 ^ x37 ;
  assign n1019 = ~n1017 & ~n1018 ;
  assign n1020 = x68 ^ x38 ;
  assign n1021 = n1019 & ~n1020 ;
  assign n1022 = n1016 & ~n1021 ;
  assign n1023 = x69 ^ x36 ;
  assign n1024 = x70 ^ x37 ;
  assign n1025 = ~n1023 & ~n1024 ;
  assign n1026 = x71 ^ x38 ;
  assign n1027 = n1025 & ~n1026 ;
  assign n1028 = n1022 & ~n1027 ;
  assign n1029 = x75 ^ x36 ;
  assign n1030 = x76 ^ x37 ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = x77 ^ x38 ;
  assign n1033 = n1031 & ~n1032 ;
  assign n1034 = n1028 & ~n1033 ;
  assign n1035 = x84 ^ x36 ;
  assign n1036 = x85 ^ x37 ;
  assign n1037 = ~n1035 & ~n1036 ;
  assign n1038 = x86 ^ x38 ;
  assign n1039 = n1037 & ~n1038 ;
  assign n1040 = n1034 & ~n1039 ;
  assign n1041 = x90 ^ x36 ;
  assign n1042 = x91 ^ x37 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = x92 ^ x38 ;
  assign n1045 = n1043 & ~n1044 ;
  assign n1046 = n1040 & ~n1045 ;
  assign n1047 = x135 ^ x36 ;
  assign n1048 = x136 ^ x37 ;
  assign n1049 = ~n1047 & ~n1048 ;
  assign n1050 = x137 ^ x38 ;
  assign n1051 = n1049 & ~n1050 ;
  assign n1052 = n1046 & ~n1051 ;
  assign n1053 = x66 ^ x39 ;
  assign n1054 = x67 ^ x40 ;
  assign n1055 = ~n1053 & ~n1054 ;
  assign n1056 = x68 ^ x41 ;
  assign n1057 = n1055 & ~n1056 ;
  assign n1058 = n1052 & ~n1057 ;
  assign n1059 = x72 ^ x39 ;
  assign n1060 = x73 ^ x40 ;
  assign n1061 = ~n1059 & ~n1060 ;
  assign n1062 = x74 ^ x41 ;
  assign n1063 = n1061 & ~n1062 ;
  assign n1064 = n1058 & ~n1063 ;
  assign n1065 = x81 ^ x39 ;
  assign n1066 = x82 ^ x40 ;
  assign n1067 = ~n1065 & ~n1066 ;
  assign n1068 = x83 ^ x41 ;
  assign n1069 = n1067 & ~n1068 ;
  assign n1070 = n1064 & ~n1069 ;
  assign n1071 = x87 ^ x39 ;
  assign n1072 = x88 ^ x40 ;
  assign n1073 = ~n1071 & ~n1072 ;
  assign n1074 = x89 ^ x41 ;
  assign n1075 = n1073 & ~n1074 ;
  assign n1076 = n1070 & ~n1075 ;
  assign n1077 = x96 ^ x39 ;
  assign n1078 = x97 ^ x40 ;
  assign n1079 = ~n1077 & ~n1078 ;
  assign n1080 = x98 ^ x41 ;
  assign n1081 = n1079 & ~n1080 ;
  assign n1082 = n1076 & ~n1081 ;
  assign n1083 = x135 ^ x39 ;
  assign n1084 = x136 ^ x40 ;
  assign n1085 = ~n1083 & ~n1084 ;
  assign n1086 = x137 ^ x41 ;
  assign n1087 = n1085 & ~n1086 ;
  assign n1088 = n1082 & ~n1087 ;
  assign n1089 = x66 ^ x42 ;
  assign n1090 = x67 ^ x43 ;
  assign n1091 = ~n1089 & ~n1090 ;
  assign n1092 = x68 ^ x44 ;
  assign n1093 = n1091 & ~n1092 ;
  assign n1094 = n1088 & ~n1093 ;
  assign n1095 = x69 ^ x42 ;
  assign n1096 = x70 ^ x43 ;
  assign n1097 = ~n1095 & ~n1096 ;
  assign n1098 = x71 ^ x44 ;
  assign n1099 = n1097 & ~n1098 ;
  assign n1100 = n1094 & ~n1099 ;
  assign n1101 = x81 ^ x42 ;
  assign n1102 = x82 ^ x43 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = x83 ^ x44 ;
  assign n1105 = n1103 & ~n1104 ;
  assign n1106 = n1100 & ~n1105 ;
  assign n1107 = x84 ^ x42 ;
  assign n1108 = x85 ^ x43 ;
  assign n1109 = ~n1107 & ~n1108 ;
  assign n1110 = x86 ^ x44 ;
  assign n1111 = n1109 & ~n1110 ;
  assign n1112 = n1106 & ~n1111 ;
  assign n1113 = x96 ^ x42 ;
  assign n1114 = x97 ^ x43 ;
  assign n1115 = ~n1113 & ~n1114 ;
  assign n1116 = x98 ^ x44 ;
  assign n1117 = n1115 & ~n1116 ;
  assign n1118 = n1112 & ~n1117 ;
  assign n1119 = x135 ^ x42 ;
  assign n1120 = x136 ^ x43 ;
  assign n1121 = ~n1119 & ~n1120 ;
  assign n1122 = x137 ^ x44 ;
  assign n1123 = n1121 & ~n1122 ;
  assign n1124 = n1118 & ~n1123 ;
  assign n1125 = x66 ^ x45 ;
  assign n1126 = x67 ^ x46 ;
  assign n1127 = ~n1125 & ~n1126 ;
  assign n1128 = x68 ^ x47 ;
  assign n1129 = n1127 & ~n1128 ;
  assign n1130 = n1124 & ~n1129 ;
  assign n1131 = x75 ^ x45 ;
  assign n1132 = x76 ^ x46 ;
  assign n1133 = ~n1131 & ~n1132 ;
  assign n1134 = x77 ^ x47 ;
  assign n1135 = n1133 & ~n1134 ;
  assign n1136 = n1130 & ~n1135 ;
  assign n1137 = x78 ^ x45 ;
  assign n1138 = x79 ^ x46 ;
  assign n1139 = ~n1137 & ~n1138 ;
  assign n1140 = x80 ^ x47 ;
  assign n1141 = n1139 & ~n1140 ;
  assign n1142 = n1136 & ~n1141 ;
  assign n1143 = x90 ^ x45 ;
  assign n1144 = x91 ^ x46 ;
  assign n1145 = ~n1143 & ~n1144 ;
  assign n1146 = x92 ^ x47 ;
  assign n1147 = n1145 & ~n1146 ;
  assign n1148 = n1142 & ~n1147 ;
  assign n1149 = x93 ^ x45 ;
  assign n1150 = x94 ^ x46 ;
  assign n1151 = ~n1149 & ~n1150 ;
  assign n1152 = x95 ^ x47 ;
  assign n1153 = n1151 & ~n1152 ;
  assign n1154 = n1148 & ~n1153 ;
  assign n1155 = x135 ^ x45 ;
  assign n1156 = x136 ^ x46 ;
  assign n1157 = ~n1155 & ~n1156 ;
  assign n1158 = x137 ^ x47 ;
  assign n1159 = n1157 & ~n1158 ;
  assign n1160 = n1154 & ~n1159 ;
  assign n1161 = x66 ^ x48 ;
  assign n1162 = x67 ^ x49 ;
  assign n1163 = ~n1161 & ~n1162 ;
  assign n1164 = x68 ^ x50 ;
  assign n1165 = n1163 & ~n1164 ;
  assign n1166 = n1160 & ~n1165 ;
  assign n1167 = x72 ^ x48 ;
  assign n1168 = x73 ^ x49 ;
  assign n1169 = ~n1167 & ~n1168 ;
  assign n1170 = x74 ^ x50 ;
  assign n1171 = n1169 & ~n1170 ;
  assign n1172 = n1166 & ~n1171 ;
  assign n1173 = x78 ^ x48 ;
  assign n1174 = x79 ^ x49 ;
  assign n1175 = ~n1173 & ~n1174 ;
  assign n1176 = x80 ^ x50 ;
  assign n1177 = n1175 & ~n1176 ;
  assign n1178 = n1172 & ~n1177 ;
  assign n1179 = x99 ^ x48 ;
  assign n1180 = x100 ^ x49 ;
  assign n1181 = ~n1179 & ~n1180 ;
  assign n1182 = x101 ^ x50 ;
  assign n1183 = n1181 & ~n1182 ;
  assign n1184 = n1178 & ~n1183 ;
  assign n1185 = x135 ^ x48 ;
  assign n1186 = x136 ^ x49 ;
  assign n1187 = ~n1185 & ~n1186 ;
  assign n1188 = x137 ^ x50 ;
  assign n1189 = n1187 & ~n1188 ;
  assign n1190 = n1184 & ~n1189 ;
  assign n1191 = x66 ^ x51 ;
  assign n1192 = x67 ^ x52 ;
  assign n1193 = ~n1191 & ~n1192 ;
  assign n1194 = x68 ^ x53 ;
  assign n1195 = n1193 & ~n1194 ;
  assign n1196 = n1190 & ~n1195 ;
  assign n1197 = x69 ^ x51 ;
  assign n1198 = x70 ^ x52 ;
  assign n1199 = ~n1197 & ~n1198 ;
  assign n1200 = x71 ^ x53 ;
  assign n1201 = n1199 & ~n1200 ;
  assign n1202 = n1196 & ~n1201 ;
  assign n1203 = x75 ^ x51 ;
  assign n1204 = x76 ^ x52 ;
  assign n1205 = ~n1203 & ~n1204 ;
  assign n1206 = x77 ^ x53 ;
  assign n1207 = n1205 & ~n1206 ;
  assign n1208 = n1202 & ~n1207 ;
  assign n1209 = x99 ^ x51 ;
  assign n1210 = x100 ^ x52 ;
  assign n1211 = ~n1209 & ~n1210 ;
  assign n1212 = x101 ^ x53 ;
  assign n1213 = n1211 & ~n1212 ;
  assign n1214 = n1208 & ~n1213 ;
  assign n1215 = x135 ^ x51 ;
  assign n1216 = x136 ^ x52 ;
  assign n1217 = ~n1215 & ~n1216 ;
  assign n1218 = x137 ^ x53 ;
  assign n1219 = n1217 & ~n1218 ;
  assign n1220 = n1214 & ~n1219 ;
  assign n1221 = x66 ^ x54 ;
  assign n1222 = x67 ^ x55 ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = x68 ^ x56 ;
  assign n1225 = n1223 & ~n1224 ;
  assign n1226 = n1220 & ~n1225 ;
  assign n1227 = x72 ^ x54 ;
  assign n1228 = x73 ^ x55 ;
  assign n1229 = ~n1227 & ~n1228 ;
  assign n1230 = x74 ^ x56 ;
  assign n1231 = n1229 & ~n1230 ;
  assign n1232 = n1226 & ~n1231 ;
  assign n1233 = x81 ^ x54 ;
  assign n1234 = x82 ^ x55 ;
  assign n1235 = ~n1233 & ~n1234 ;
  assign n1236 = x83 ^ x56 ;
  assign n1237 = n1235 & ~n1236 ;
  assign n1238 = n1232 & ~n1237 ;
  assign n1239 = x99 ^ x54 ;
  assign n1240 = x100 ^ x55 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = x101 ^ x56 ;
  assign n1243 = n1241 & ~n1242 ;
  assign n1244 = n1238 & ~n1243 ;
  assign n1245 = x135 ^ x54 ;
  assign n1246 = x136 ^ x55 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = x137 ^ x56 ;
  assign n1249 = n1247 & ~n1248 ;
  assign n1250 = n1244 & ~n1249 ;
  assign n1251 = x66 ^ x57 ;
  assign n1252 = x67 ^ x58 ;
  assign n1253 = ~n1251 & ~n1252 ;
  assign n1254 = x68 ^ x59 ;
  assign n1255 = n1253 & ~n1254 ;
  assign n1256 = n1250 & ~n1255 ;
  assign n1257 = x69 ^ x57 ;
  assign n1258 = x70 ^ x58 ;
  assign n1259 = ~n1257 & ~n1258 ;
  assign n1260 = x71 ^ x59 ;
  assign n1261 = n1259 & ~n1260 ;
  assign n1262 = n1256 & ~n1261 ;
  assign n1263 = x81 ^ x57 ;
  assign n1264 = x82 ^ x58 ;
  assign n1265 = ~n1263 & ~n1264 ;
  assign n1266 = x83 ^ x59 ;
  assign n1267 = n1265 & ~n1266 ;
  assign n1268 = n1262 & ~n1267 ;
  assign n1269 = x99 ^ x57 ;
  assign n1270 = x100 ^ x58 ;
  assign n1271 = ~n1269 & ~n1270 ;
  assign n1272 = x101 ^ x59 ;
  assign n1273 = n1271 & ~n1272 ;
  assign n1274 = n1268 & ~n1273 ;
  assign n1275 = x135 ^ x57 ;
  assign n1276 = x136 ^ x58 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1278 = x137 ^ x59 ;
  assign n1279 = n1277 & ~n1278 ;
  assign n1280 = n1274 & ~n1279 ;
  assign n1281 = x66 ^ x60 ;
  assign n1282 = x67 ^ x61 ;
  assign n1283 = ~n1281 & ~n1282 ;
  assign n1284 = x68 ^ x62 ;
  assign n1285 = n1283 & ~n1284 ;
  assign n1286 = n1280 & ~n1285 ;
  assign n1287 = x75 ^ x60 ;
  assign n1288 = x76 ^ x61 ;
  assign n1289 = ~n1287 & ~n1288 ;
  assign n1290 = x77 ^ x62 ;
  assign n1291 = n1289 & ~n1290 ;
  assign n1292 = n1286 & ~n1291 ;
  assign n1293 = x78 ^ x60 ;
  assign n1294 = x79 ^ x61 ;
  assign n1295 = ~n1293 & ~n1294 ;
  assign n1296 = x80 ^ x62 ;
  assign n1297 = n1295 & ~n1296 ;
  assign n1298 = n1292 & ~n1297 ;
  assign n1299 = x99 ^ x60 ;
  assign n1300 = x100 ^ x61 ;
  assign n1301 = ~n1299 & ~n1300 ;
  assign n1302 = x101 ^ x62 ;
  assign n1303 = n1301 & ~n1302 ;
  assign n1304 = n1298 & ~n1303 ;
  assign n1305 = x135 ^ x60 ;
  assign n1306 = x136 ^ x61 ;
  assign n1307 = ~n1305 & ~n1306 ;
  assign n1308 = x137 ^ x62 ;
  assign n1309 = n1307 & ~n1308 ;
  assign n1310 = n1304 & ~n1309 ;
  assign n1311 = x66 ^ x63 ;
  assign n1312 = x67 ^ x64 ;
  assign n1313 = ~n1311 & ~n1312 ;
  assign n1314 = x68 ^ x65 ;
  assign n1315 = n1313 & ~n1314 ;
  assign n1316 = n1310 & ~n1315 ;
  assign n1317 = x84 ^ x63 ;
  assign n1318 = x85 ^ x64 ;
  assign n1319 = ~n1317 & ~n1318 ;
  assign n1320 = x86 ^ x65 ;
  assign n1321 = n1319 & ~n1320 ;
  assign n1322 = n1316 & ~n1321 ;
  assign n1323 = x87 ^ x63 ;
  assign n1324 = x88 ^ x64 ;
  assign n1325 = ~n1323 & ~n1324 ;
  assign n1326 = x89 ^ x65 ;
  assign n1327 = n1325 & ~n1326 ;
  assign n1328 = n1322 & ~n1327 ;
  assign n1329 = x90 ^ x63 ;
  assign n1330 = x91 ^ x64 ;
  assign n1331 = ~n1329 & ~n1330 ;
  assign n1332 = x92 ^ x65 ;
  assign n1333 = n1331 & ~n1332 ;
  assign n1334 = n1328 & ~n1333 ;
  assign n1335 = x93 ^ x63 ;
  assign n1336 = x94 ^ x64 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = x95 ^ x65 ;
  assign n1339 = n1337 & ~n1338 ;
  assign n1340 = n1334 & ~n1339 ;
  assign n1341 = x96 ^ x63 ;
  assign n1342 = x97 ^ x64 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = x98 ^ x65 ;
  assign n1345 = n1343 & ~n1344 ;
  assign n1346 = n1340 & ~n1345 ;
  assign n1347 = x135 ^ x63 ;
  assign n1348 = x136 ^ x64 ;
  assign n1349 = ~n1347 & ~n1348 ;
  assign n1350 = x137 ^ x65 ;
  assign n1351 = n1349 & ~n1350 ;
  assign n1352 = n1346 & ~n1351 ;
  assign n1353 = x102 ^ x66 ;
  assign n1354 = x103 ^ x67 ;
  assign n1355 = ~n1353 & ~n1354 ;
  assign n1356 = x104 ^ x68 ;
  assign n1357 = n1355 & ~n1356 ;
  assign n1358 = n1352 & ~n1357 ;
  assign n1359 = x105 ^ x66 ;
  assign n1360 = x106 ^ x67 ;
  assign n1361 = ~n1359 & ~n1360 ;
  assign n1362 = x107 ^ x68 ;
  assign n1363 = n1361 & ~n1362 ;
  assign n1364 = n1358 & ~n1363 ;
  assign n1365 = x108 ^ x66 ;
  assign n1366 = x109 ^ x67 ;
  assign n1367 = ~n1365 & ~n1366 ;
  assign n1368 = x110 ^ x68 ;
  assign n1369 = n1367 & ~n1368 ;
  assign n1370 = n1364 & ~n1369 ;
  assign n1371 = x111 ^ x66 ;
  assign n1372 = x112 ^ x67 ;
  assign n1373 = ~n1371 & ~n1372 ;
  assign n1374 = x113 ^ x68 ;
  assign n1375 = n1373 & ~n1374 ;
  assign n1376 = n1370 & ~n1375 ;
  assign n1377 = x114 ^ x66 ;
  assign n1378 = x115 ^ x67 ;
  assign n1379 = ~n1377 & ~n1378 ;
  assign n1380 = x116 ^ x68 ;
  assign n1381 = n1379 & ~n1380 ;
  assign n1382 = n1376 & ~n1381 ;
  assign n1383 = x117 ^ x66 ;
  assign n1384 = x118 ^ x67 ;
  assign n1385 = ~n1383 & ~n1384 ;
  assign n1386 = x119 ^ x68 ;
  assign n1387 = n1385 & ~n1386 ;
  assign n1388 = n1382 & ~n1387 ;
  assign n1389 = x120 ^ x66 ;
  assign n1390 = x121 ^ x67 ;
  assign n1391 = ~n1389 & ~n1390 ;
  assign n1392 = x122 ^ x68 ;
  assign n1393 = n1391 & ~n1392 ;
  assign n1394 = n1388 & ~n1393 ;
  assign n1395 = x123 ^ x66 ;
  assign n1396 = x124 ^ x67 ;
  assign n1397 = ~n1395 & ~n1396 ;
  assign n1398 = x125 ^ x68 ;
  assign n1399 = n1397 & ~n1398 ;
  assign n1400 = n1394 & ~n1399 ;
  assign n1401 = x126 ^ x66 ;
  assign n1402 = x127 ^ x67 ;
  assign n1403 = ~n1401 & ~n1402 ;
  assign n1404 = x128 ^ x68 ;
  assign n1405 = n1403 & ~n1404 ;
  assign n1406 = n1400 & ~n1405 ;
  assign n1407 = x129 ^ x66 ;
  assign n1408 = x130 ^ x67 ;
  assign n1409 = ~n1407 & ~n1408 ;
  assign n1410 = x131 ^ x68 ;
  assign n1411 = n1409 & ~n1410 ;
  assign n1412 = n1406 & ~n1411 ;
  assign n1413 = x132 ^ x66 ;
  assign n1414 = x133 ^ x67 ;
  assign n1415 = ~n1413 & ~n1414 ;
  assign n1416 = x134 ^ x68 ;
  assign n1417 = n1415 & ~n1416 ;
  assign n1418 = n1412 & ~n1417 ;
  assign n1419 = x138 ^ x69 ;
  assign n1420 = x139 ^ x70 ;
  assign n1421 = ~n1419 & ~n1420 ;
  assign n1422 = x140 ^ x71 ;
  assign n1423 = n1421 & ~n1422 ;
  assign n1424 = n1418 & ~n1423 ;
  assign n1425 = x138 ^ x72 ;
  assign n1426 = x139 ^ x73 ;
  assign n1427 = ~n1425 & ~n1426 ;
  assign n1428 = x140 ^ x74 ;
  assign n1429 = n1427 & ~n1428 ;
  assign n1430 = n1424 & ~n1429 ;
  assign n1431 = x138 ^ x75 ;
  assign n1432 = x139 ^ x76 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = x140 ^ x77 ;
  assign n1435 = n1433 & ~n1434 ;
  assign n1436 = n1430 & ~n1435 ;
  assign n1437 = x138 ^ x78 ;
  assign n1438 = x139 ^ x79 ;
  assign n1439 = ~n1437 & ~n1438 ;
  assign n1440 = x140 ^ x80 ;
  assign n1441 = n1439 & ~n1440 ;
  assign n1442 = n1436 & ~n1441 ;
  assign n1443 = x138 ^ x81 ;
  assign n1444 = x139 ^ x82 ;
  assign n1445 = ~n1443 & ~n1444 ;
  assign n1446 = x140 ^ x83 ;
  assign n1447 = n1445 & ~n1446 ;
  assign n1448 = n1442 & ~n1447 ;
  assign n1449 = x138 ^ x84 ;
  assign n1450 = x139 ^ x85 ;
  assign n1451 = ~n1449 & ~n1450 ;
  assign n1452 = x140 ^ x86 ;
  assign n1453 = n1451 & ~n1452 ;
  assign n1454 = n1448 & ~n1453 ;
  assign n1455 = x138 ^ x87 ;
  assign n1456 = x139 ^ x88 ;
  assign n1457 = ~n1455 & ~n1456 ;
  assign n1458 = x140 ^ x89 ;
  assign n1459 = n1457 & ~n1458 ;
  assign n1460 = n1454 & ~n1459 ;
  assign n1461 = x138 ^ x90 ;
  assign n1462 = x139 ^ x91 ;
  assign n1463 = ~n1461 & ~n1462 ;
  assign n1464 = x140 ^ x92 ;
  assign n1465 = n1463 & ~n1464 ;
  assign n1466 = n1460 & ~n1465 ;
  assign n1467 = x138 ^ x93 ;
  assign n1468 = x139 ^ x94 ;
  assign n1469 = ~n1467 & ~n1468 ;
  assign n1470 = x140 ^ x95 ;
  assign n1471 = n1469 & ~n1470 ;
  assign n1472 = n1466 & ~n1471 ;
  assign n1473 = x138 ^ x96 ;
  assign n1474 = x139 ^ x97 ;
  assign n1475 = ~n1473 & ~n1474 ;
  assign n1476 = x140 ^ x98 ;
  assign n1477 = n1475 & ~n1476 ;
  assign n1478 = n1472 & ~n1477 ;
  assign n1479 = x138 ^ x99 ;
  assign n1480 = x139 ^ x100 ;
  assign n1481 = ~n1479 & ~n1480 ;
  assign n1482 = x140 ^ x101 ;
  assign n1483 = n1481 & ~n1482 ;
  assign n1484 = n1478 & ~n1483 ;
  assign n1485 = x138 ^ x102 ;
  assign n1486 = x139 ^ x103 ;
  assign n1487 = ~n1485 & ~n1486 ;
  assign n1488 = x140 ^ x104 ;
  assign n1489 = n1487 & ~n1488 ;
  assign n1490 = n1484 & ~n1489 ;
  assign n1491 = x138 ^ x105 ;
  assign n1492 = x139 ^ x106 ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1494 = x140 ^ x107 ;
  assign n1495 = n1493 & ~n1494 ;
  assign n1496 = n1490 & ~n1495 ;
  assign n1497 = x138 ^ x108 ;
  assign n1498 = x139 ^ x109 ;
  assign n1499 = ~n1497 & ~n1498 ;
  assign n1500 = x140 ^ x110 ;
  assign n1501 = n1499 & ~n1500 ;
  assign n1502 = n1496 & ~n1501 ;
  assign n1503 = x138 ^ x111 ;
  assign n1504 = x139 ^ x112 ;
  assign n1505 = ~n1503 & ~n1504 ;
  assign n1506 = x140 ^ x113 ;
  assign n1507 = n1505 & ~n1506 ;
  assign n1508 = n1502 & ~n1507 ;
  assign n1509 = x138 ^ x114 ;
  assign n1510 = x139 ^ x115 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = x140 ^ x116 ;
  assign n1513 = n1511 & ~n1512 ;
  assign n1514 = n1508 & ~n1513 ;
  assign n1515 = x138 ^ x117 ;
  assign n1516 = x139 ^ x118 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1518 = x140 ^ x119 ;
  assign n1519 = n1517 & ~n1518 ;
  assign n1520 = n1514 & ~n1519 ;
  assign n1521 = x138 ^ x120 ;
  assign n1522 = x139 ^ x121 ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = x140 ^ x122 ;
  assign n1525 = n1523 & ~n1524 ;
  assign n1526 = n1520 & ~n1525 ;
  assign n1527 = x138 ^ x123 ;
  assign n1528 = x139 ^ x124 ;
  assign n1529 = ~n1527 & ~n1528 ;
  assign n1530 = x140 ^ x125 ;
  assign n1531 = n1529 & ~n1530 ;
  assign n1532 = n1526 & ~n1531 ;
  assign n1533 = x138 ^ x126 ;
  assign n1534 = x139 ^ x127 ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1536 = x140 ^ x128 ;
  assign n1537 = n1535 & ~n1536 ;
  assign n1538 = n1532 & ~n1537 ;
  assign n1539 = x138 ^ x129 ;
  assign n1540 = x139 ^ x130 ;
  assign n1541 = ~n1539 & ~n1540 ;
  assign n1542 = x140 ^ x131 ;
  assign n1543 = n1541 & ~n1542 ;
  assign n1544 = n1538 & ~n1543 ;
  assign n1545 = x138 ^ x132 ;
  assign n1546 = x139 ^ x133 ;
  assign n1547 = ~n1545 & ~n1546 ;
  assign n1548 = x140 ^ x134 ;
  assign n1549 = n1547 & ~n1548 ;
  assign n1550 = n1544 & ~n1549 ;
  assign n1551 = x138 ^ x135 ;
  assign n1552 = x139 ^ x136 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = x140 ^ x137 ;
  assign n1555 = n1553 & ~n1554 ;
  assign n1556 = n1550 & ~n1555 ;
  assign y0 = n1556 ;
endmodule
