module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n13 = x2 ^ x0 ;
  assign n14 = x3 ^ x1 ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = x4 ^ x2 ;
  assign n17 = x5 ^ x3 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = ~n15 & ~n18 ;
  assign n20 = x10 ^ x2 ;
  assign n21 = x11 ^ x3 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = n19 & ~n22 ;
  assign n24 = x6 ^ x4 ;
  assign n25 = x7 ^ x5 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = n23 & ~n26 ;
  assign n28 = x8 ^ x6 ;
  assign n29 = x9 ^ x7 ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = n27 & ~n30 ;
  assign y0 = n31 ;
endmodule
