module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n13 = x2 ^ x0 ;
  assign n14 = x3 ^ x1 ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = x4 ^ x2 ;
  assign n17 = x5 ^ x3 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = x10 ^ x2 ;
  assign n20 = x11 ^ x3 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = x6 ^ x4 ;
  assign n23 = x7 ^ x5 ;
  assign n24 = ~n22 & ~n23 ;
  assign n25 = x8 ^ x6 ;
  assign n26 = x9 ^ x7 ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = ~n15 & ~n18 ;
  assign n29 = n28 & ~n21 ;
  assign n30 = n29 & ~n24 ;
  assign y0 = n30 & ~n27 ;
endmodule
