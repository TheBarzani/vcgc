module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 ;
  assign n61 = x2 ^ x0 ;
  assign n62 = x3 ^ x1 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = x6 ^ x0 ;
  assign n65 = x7 ^ x1 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = ~n63 & ~n66 ;
  assign n68 = x20 ^ x0 ;
  assign n69 = x21 ^ x1 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = n67 & ~n70 ;
  assign n72 = x24 ^ x0 ;
  assign n73 = x25 ^ x1 ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = n71 & ~n74 ;
  assign n76 = x4 ^ x2 ;
  assign n77 = x5 ^ x3 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = n75 & ~n78 ;
  assign n80 = x18 ^ x2 ;
  assign n81 = x19 ^ x3 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = n79 & ~n82 ;
  assign n84 = x22 ^ x2 ;
  assign n85 = x23 ^ x3 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n83 & ~n86 ;
  assign n88 = x10 ^ x4 ;
  assign n89 = x11 ^ x5 ;
  assign n90 = ~n88 & ~n89 ;
  assign n91 = n87 & ~n90 ;
  assign n92 = x14 ^ x4 ;
  assign n93 = x15 ^ x5 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = n91 & ~n94 ;
  assign n96 = x20 ^ x4 ;
  assign n97 = x21 ^ x5 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = n95 & ~n98 ;
  assign n100 = x28 ^ x4 ;
  assign n101 = x29 ^ x5 ;
  assign n102 = ~n100 & ~n101 ;
  assign n103 = n99 & ~n102 ;
  assign n104 = x32 ^ x4 ;
  assign n105 = x33 ^ x5 ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = n103 & ~n106 ;
  assign n108 = x8 ^ x6 ;
  assign n109 = x9 ^ x7 ;
  assign n110 = ~n108 & ~n109 ;
  assign n111 = n107 & ~n110 ;
  assign n112 = x14 ^ x6 ;
  assign n113 = x15 ^ x7 ;
  assign n114 = ~n112 & ~n113 ;
  assign n115 = n111 & ~n114 ;
  assign n116 = x18 ^ x6 ;
  assign n117 = x19 ^ x7 ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = n115 & ~n118 ;
  assign n120 = x26 ^ x6 ;
  assign n121 = x27 ^ x7 ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = n119 & ~n122 ;
  assign n124 = x32 ^ x6 ;
  assign n125 = x33 ^ x7 ;
  assign n126 = ~n124 & ~n125 ;
  assign n127 = n123 & ~n126 ;
  assign n128 = x12 ^ x8 ;
  assign n129 = x13 ^ x9 ;
  assign n130 = ~n128 & ~n129 ;
  assign n131 = n127 & ~n130 ;
  assign n132 = x16 ^ x8 ;
  assign n133 = x17 ^ x9 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = n131 & ~n134 ;
  assign n136 = x24 ^ x8 ;
  assign n137 = x25 ^ x9 ;
  assign n138 = ~n136 & ~n137 ;
  assign n139 = n135 & ~n138 ;
  assign n140 = x30 ^ x8 ;
  assign n141 = x31 ^ x9 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n139 & ~n142 ;
  assign n144 = x34 ^ x8 ;
  assign n145 = x35 ^ x9 ;
  assign n146 = ~n144 & ~n145 ;
  assign n147 = n143 & ~n146 ;
  assign n148 = x12 ^ x10 ;
  assign n149 = x13 ^ x11 ;
  assign n150 = ~n148 & ~n149 ;
  assign n151 = n147 & ~n150 ;
  assign n152 = x16 ^ x10 ;
  assign n153 = x17 ^ x11 ;
  assign n154 = ~n152 & ~n153 ;
  assign n155 = n151 & ~n154 ;
  assign n156 = x22 ^ x10 ;
  assign n157 = x23 ^ x11 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = n155 & ~n158 ;
  assign n160 = x30 ^ x10 ;
  assign n161 = x31 ^ x11 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = n159 & ~n162 ;
  assign n164 = x34 ^ x10 ;
  assign n165 = x35 ^ x11 ;
  assign n166 = ~n164 & ~n165 ;
  assign n167 = n163 & ~n166 ;
  assign n168 = x14 ^ x12 ;
  assign n169 = x15 ^ x13 ;
  assign n170 = ~n168 & ~n169 ;
  assign n171 = n167 & ~n170 ;
  assign n172 = x16 ^ x12 ;
  assign n173 = x17 ^ x13 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = n171 & ~n174 ;
  assign n176 = x26 ^ x12 ;
  assign n177 = x27 ^ x13 ;
  assign n178 = ~n176 & ~n177 ;
  assign n179 = n175 & ~n178 ;
  assign n180 = x28 ^ x12 ;
  assign n181 = x29 ^ x13 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = n179 & ~n182 ;
  assign n184 = x32 ^ x12 ;
  assign n185 = x33 ^ x13 ;
  assign n186 = ~n184 & ~n185 ;
  assign n187 = n183 & ~n186 ;
  assign n188 = x34 ^ x12 ;
  assign n189 = x35 ^ x13 ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = n187 & ~n190 ;
  assign n192 = x16 ^ x14 ;
  assign n193 = x17 ^ x15 ;
  assign n194 = ~n192 & ~n193 ;
  assign n195 = n191 & ~n194 ;
  assign n196 = x22 ^ x14 ;
  assign n197 = x23 ^ x15 ;
  assign n198 = ~n196 & ~n197 ;
  assign n199 = n195 & ~n198 ;
  assign n200 = x24 ^ x14 ;
  assign n201 = x25 ^ x15 ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = n199 & ~n202 ;
  assign n204 = x30 ^ x14 ;
  assign n205 = x31 ^ x15 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = n203 & ~n206 ;
  assign n208 = x34 ^ x14 ;
  assign n209 = x35 ^ x15 ;
  assign n210 = ~n208 & ~n209 ;
  assign n211 = n207 & ~n210 ;
  assign n212 = x26 ^ x16 ;
  assign n213 = x27 ^ x17 ;
  assign n214 = ~n212 & ~n213 ;
  assign n215 = n211 & ~n214 ;
  assign n216 = x28 ^ x16 ;
  assign n217 = x29 ^ x17 ;
  assign n218 = ~n216 & ~n217 ;
  assign n219 = n215 & ~n218 ;
  assign n220 = x30 ^ x16 ;
  assign n221 = x31 ^ x17 ;
  assign n222 = ~n220 & ~n221 ;
  assign n223 = n219 & ~n222 ;
  assign n224 = x32 ^ x16 ;
  assign n225 = x33 ^ x17 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = n223 & ~n226 ;
  assign n228 = x38 ^ x18 ;
  assign n229 = x39 ^ x19 ;
  assign n230 = ~n228 & ~n229 ;
  assign n231 = n227 & ~n230 ;
  assign n232 = x42 ^ x18 ;
  assign n233 = x43 ^ x19 ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = n231 & ~n234 ;
  assign n236 = x56 ^ x18 ;
  assign n237 = x57 ^ x19 ;
  assign n238 = ~n236 & ~n237 ;
  assign n239 = n235 & ~n238 ;
  assign n240 = x36 ^ x20 ;
  assign n241 = x37 ^ x21 ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = n239 & ~n242 ;
  assign n244 = x40 ^ x20 ;
  assign n245 = x41 ^ x21 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = n243 & ~n246 ;
  assign n248 = x56 ^ x20 ;
  assign n249 = x57 ^ x21 ;
  assign n250 = ~n248 & ~n249 ;
  assign n251 = n247 & ~n250 ;
  assign n252 = x38 ^ x22 ;
  assign n253 = x39 ^ x23 ;
  assign n254 = ~n252 & ~n253 ;
  assign n255 = n251 & ~n254 ;
  assign n256 = x46 ^ x22 ;
  assign n257 = x47 ^ x23 ;
  assign n258 = ~n256 & ~n257 ;
  assign n259 = n255 & ~n258 ;
  assign n260 = x50 ^ x22 ;
  assign n261 = x51 ^ x23 ;
  assign n262 = ~n260 & ~n261 ;
  assign n263 = n259 & ~n262 ;
  assign n264 = x56 ^ x22 ;
  assign n265 = x57 ^ x23 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n263 & ~n266 ;
  assign n268 = x36 ^ x24 ;
  assign n269 = x37 ^ x25 ;
  assign n270 = ~n268 & ~n269 ;
  assign n271 = n267 & ~n270 ;
  assign n272 = x44 ^ x24 ;
  assign n273 = x45 ^ x25 ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = n271 & ~n274 ;
  assign n276 = x50 ^ x24 ;
  assign n277 = x51 ^ x25 ;
  assign n278 = ~n276 & ~n277 ;
  assign n279 = n275 & ~n278 ;
  assign n280 = x56 ^ x24 ;
  assign n281 = x57 ^ x25 ;
  assign n282 = ~n280 & ~n281 ;
  assign n283 = n279 & ~n282 ;
  assign n284 = x42 ^ x26 ;
  assign n285 = x43 ^ x27 ;
  assign n286 = ~n284 & ~n285 ;
  assign n287 = n283 & ~n286 ;
  assign n288 = x48 ^ x26 ;
  assign n289 = x49 ^ x27 ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = n287 & ~n290 ;
  assign n292 = x52 ^ x26 ;
  assign n293 = x53 ^ x27 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = n291 & ~n294 ;
  assign n296 = x56 ^ x26 ;
  assign n297 = x57 ^ x27 ;
  assign n298 = ~n296 & ~n297 ;
  assign n299 = n295 & ~n298 ;
  assign n300 = x40 ^ x28 ;
  assign n301 = x41 ^ x29 ;
  assign n302 = ~n300 & ~n301 ;
  assign n303 = n299 & ~n302 ;
  assign n304 = x48 ^ x28 ;
  assign n305 = x49 ^ x29 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = n303 & ~n306 ;
  assign n308 = x52 ^ x28 ;
  assign n309 = x53 ^ x29 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = n307 & ~n310 ;
  assign n312 = x56 ^ x28 ;
  assign n313 = x57 ^ x29 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = n311 & ~n314 ;
  assign n316 = x44 ^ x30 ;
  assign n317 = x45 ^ x31 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = n315 & ~n318 ;
  assign n320 = x46 ^ x30 ;
  assign n321 = x47 ^ x31 ;
  assign n322 = ~n320 & ~n321 ;
  assign n323 = n319 & ~n322 ;
  assign n324 = x50 ^ x30 ;
  assign n325 = x51 ^ x31 ;
  assign n326 = ~n324 & ~n325 ;
  assign n327 = n323 & ~n326 ;
  assign n328 = x52 ^ x30 ;
  assign n329 = x53 ^ x31 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = n327 & ~n330 ;
  assign n332 = x56 ^ x30 ;
  assign n333 = x57 ^ x31 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = n331 & ~n334 ;
  assign n336 = x40 ^ x32 ;
  assign n337 = x41 ^ x33 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = n335 & ~n338 ;
  assign n340 = x42 ^ x32 ;
  assign n341 = x43 ^ x33 ;
  assign n342 = ~n340 & ~n341 ;
  assign n343 = n339 & ~n342 ;
  assign n344 = x48 ^ x32 ;
  assign n345 = x49 ^ x33 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = n343 & ~n346 ;
  assign n348 = x52 ^ x32 ;
  assign n349 = x53 ^ x33 ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = n347 & ~n350 ;
  assign n352 = x56 ^ x32 ;
  assign n353 = x57 ^ x33 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = n351 & ~n354 ;
  assign n356 = x44 ^ x34 ;
  assign n357 = x45 ^ x35 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = n355 & ~n358 ;
  assign n360 = x46 ^ x34 ;
  assign n361 = x47 ^ x35 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = n359 & ~n362 ;
  assign n364 = x48 ^ x34 ;
  assign n365 = x49 ^ x35 ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = n363 & ~n366 ;
  assign n368 = x50 ^ x34 ;
  assign n369 = x51 ^ x35 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = n367 & ~n370 ;
  assign n372 = x56 ^ x34 ;
  assign n373 = x57 ^ x35 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = n371 & ~n374 ;
  assign n376 = x54 ^ x36 ;
  assign n377 = x55 ^ x37 ;
  assign n378 = ~n376 & ~n377 ;
  assign n379 = n375 & ~n378 ;
  assign n380 = x58 ^ x36 ;
  assign n381 = x59 ^ x37 ;
  assign n382 = ~n380 & ~n381 ;
  assign n383 = n379 & ~n382 ;
  assign n384 = x54 ^ x38 ;
  assign n385 = x55 ^ x39 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = n383 & ~n386 ;
  assign n388 = x58 ^ x38 ;
  assign n389 = x59 ^ x39 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = n387 & ~n390 ;
  assign n392 = x54 ^ x40 ;
  assign n393 = x55 ^ x41 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = n391 & ~n394 ;
  assign n396 = x58 ^ x40 ;
  assign n397 = x59 ^ x41 ;
  assign n398 = ~n396 & ~n397 ;
  assign n399 = n395 & ~n398 ;
  assign n400 = x54 ^ x42 ;
  assign n401 = x55 ^ x43 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = n399 & ~n402 ;
  assign n404 = x58 ^ x42 ;
  assign n405 = x59 ^ x43 ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = n403 & ~n406 ;
  assign n408 = x54 ^ x44 ;
  assign n409 = x55 ^ x45 ;
  assign n410 = ~n408 & ~n409 ;
  assign n411 = n407 & ~n410 ;
  assign n412 = x58 ^ x44 ;
  assign n413 = x59 ^ x45 ;
  assign n414 = ~n412 & ~n413 ;
  assign n415 = n411 & ~n414 ;
  assign n416 = x54 ^ x46 ;
  assign n417 = x55 ^ x47 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = n415 & ~n418 ;
  assign n420 = x58 ^ x46 ;
  assign n421 = x59 ^ x47 ;
  assign n422 = ~n420 & ~n421 ;
  assign n423 = n419 & ~n422 ;
  assign n424 = x54 ^ x48 ;
  assign n425 = x55 ^ x49 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = n423 & ~n426 ;
  assign n428 = x58 ^ x48 ;
  assign n429 = x59 ^ x49 ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = n427 & ~n430 ;
  assign n432 = x54 ^ x50 ;
  assign n433 = x55 ^ x51 ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = n431 & ~n434 ;
  assign n436 = x58 ^ x50 ;
  assign n437 = x59 ^ x51 ;
  assign n438 = ~n436 & ~n437 ;
  assign n439 = n435 & ~n438 ;
  assign n440 = x54 ^ x52 ;
  assign n441 = x55 ^ x53 ;
  assign n442 = ~n440 & ~n441 ;
  assign n443 = n439 & ~n442 ;
  assign n444 = x58 ^ x52 ;
  assign n445 = x59 ^ x53 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = n443 & ~n446 ;
  assign n448 = x56 ^ x54 ;
  assign n449 = x57 ^ x55 ;
  assign n450 = ~n448 & ~n449 ;
  assign n451 = n447 & ~n450 ;
  assign n452 = x58 ^ x54 ;
  assign n453 = x59 ^ x55 ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = n451 & ~n454 ;
  assign n456 = x58 ^ x56 ;
  assign n457 = x59 ^ x57 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = n455 & ~n458 ;
  assign y0 = n459 ;
endmodule
