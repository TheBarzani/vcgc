module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 ;
  output y0 ;
  wire n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 ;
  assign n70 = x3 ^ x0 ;
  assign n71 = x4 ^ x1 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = x5 ^ x2 ;
  assign n74 = n72 & ~n73 ;
  assign n75 = x9 ^ x0 ;
  assign n76 = x10 ^ x1 ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = x11 ^ x2 ;
  assign n79 = n77 & ~n78 ;
  assign n80 = ~n74 & ~n79 ;
  assign n81 = x18 ^ x0 ;
  assign n82 = x19 ^ x1 ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = x20 ^ x2 ;
  assign n85 = n83 & ~n84 ;
  assign n86 = n80 & ~n85 ;
  assign n87 = x24 ^ x0 ;
  assign n88 = x25 ^ x1 ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = x26 ^ x2 ;
  assign n91 = n89 & ~n90 ;
  assign n92 = n86 & ~n91 ;
  assign n93 = x36 ^ x0 ;
  assign n94 = x37 ^ x1 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = x38 ^ x2 ;
  assign n97 = n95 & ~n96 ;
  assign n98 = n92 & ~n97 ;
  assign n99 = x42 ^ x0 ;
  assign n100 = x43 ^ x1 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = x44 ^ x2 ;
  assign n103 = n101 & ~n102 ;
  assign n104 = n98 & ~n103 ;
  assign n105 = x51 ^ x0 ;
  assign n106 = x52 ^ x1 ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = x53 ^ x2 ;
  assign n109 = n107 & ~n108 ;
  assign n110 = n104 & ~n109 ;
  assign n111 = x57 ^ x0 ;
  assign n112 = x58 ^ x1 ;
  assign n113 = ~n111 & ~n112 ;
  assign n114 = x59 ^ x2 ;
  assign n115 = n113 & ~n114 ;
  assign n116 = n110 & ~n115 ;
  assign n117 = x6 ^ x3 ;
  assign n118 = x7 ^ x4 ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = x8 ^ x5 ;
  assign n121 = n119 & ~n120 ;
  assign n122 = n116 & ~n121 ;
  assign n123 = x15 ^ x3 ;
  assign n124 = x16 ^ x4 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = x17 ^ x5 ;
  assign n127 = n125 & ~n126 ;
  assign n128 = n122 & ~n127 ;
  assign n129 = x21 ^ x3 ;
  assign n130 = x22 ^ x4 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = x23 ^ x5 ;
  assign n133 = n131 & ~n132 ;
  assign n134 = n128 & ~n133 ;
  assign n135 = x33 ^ x3 ;
  assign n136 = x34 ^ x4 ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = x35 ^ x5 ;
  assign n139 = n137 & ~n138 ;
  assign n140 = n134 & ~n139 ;
  assign n141 = x39 ^ x3 ;
  assign n142 = x40 ^ x4 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = x41 ^ x5 ;
  assign n145 = n143 & ~n144 ;
  assign n146 = n140 & ~n145 ;
  assign n147 = x48 ^ x3 ;
  assign n148 = x49 ^ x4 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = x50 ^ x5 ;
  assign n151 = n149 & ~n150 ;
  assign n152 = n146 & ~n151 ;
  assign n153 = x54 ^ x3 ;
  assign n154 = x55 ^ x4 ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = x56 ^ x5 ;
  assign n157 = n155 & ~n156 ;
  assign n158 = n152 & ~n157 ;
  assign n159 = x12 ^ x6 ;
  assign n160 = x13 ^ x7 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = x14 ^ x8 ;
  assign n163 = n161 & ~n162 ;
  assign n164 = n158 & ~n163 ;
  assign n165 = x18 ^ x6 ;
  assign n166 = x19 ^ x7 ;
  assign n167 = ~n165 & ~n166 ;
  assign n168 = x20 ^ x8 ;
  assign n169 = n167 & ~n168 ;
  assign n170 = n164 & ~n169 ;
  assign n171 = x27 ^ x6 ;
  assign n172 = x28 ^ x7 ;
  assign n173 = ~n171 & ~n172 ;
  assign n174 = x29 ^ x8 ;
  assign n175 = n173 & ~n174 ;
  assign n176 = n170 & ~n175 ;
  assign n177 = x36 ^ x6 ;
  assign n178 = x37 ^ x7 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = x38 ^ x8 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n176 & ~n181 ;
  assign n183 = x45 ^ x6 ;
  assign n184 = x46 ^ x7 ;
  assign n185 = ~n183 & ~n184 ;
  assign n186 = x47 ^ x8 ;
  assign n187 = n185 & ~n186 ;
  assign n188 = n182 & ~n187 ;
  assign n189 = x51 ^ x6 ;
  assign n190 = x52 ^ x7 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = x53 ^ x8 ;
  assign n193 = n191 & ~n192 ;
  assign n194 = n188 & ~n193 ;
  assign n195 = x60 ^ x6 ;
  assign n196 = x61 ^ x7 ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = x62 ^ x8 ;
  assign n199 = n197 & ~n198 ;
  assign n200 = n194 & ~n199 ;
  assign n201 = x12 ^ x9 ;
  assign n202 = x13 ^ x10 ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = x14 ^ x11 ;
  assign n205 = n203 & ~n204 ;
  assign n206 = n200 & ~n205 ;
  assign n207 = x15 ^ x9 ;
  assign n208 = x16 ^ x10 ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = x17 ^ x11 ;
  assign n211 = n209 & ~n210 ;
  assign n212 = n206 & ~n211 ;
  assign n213 = x27 ^ x9 ;
  assign n214 = x28 ^ x10 ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = x29 ^ x11 ;
  assign n217 = n215 & ~n216 ;
  assign n218 = n212 & ~n217 ;
  assign n219 = x33 ^ x9 ;
  assign n220 = x34 ^ x10 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = x35 ^ x11 ;
  assign n223 = n221 & ~n222 ;
  assign n224 = n218 & ~n223 ;
  assign n225 = x45 ^ x9 ;
  assign n226 = x46 ^ x10 ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = x47 ^ x11 ;
  assign n229 = n227 & ~n228 ;
  assign n230 = n224 & ~n229 ;
  assign n231 = x48 ^ x9 ;
  assign n232 = x49 ^ x10 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = x50 ^ x11 ;
  assign n235 = n233 & ~n234 ;
  assign n236 = n230 & ~n235 ;
  assign n237 = x60 ^ x9 ;
  assign n238 = x61 ^ x10 ;
  assign n239 = ~n237 & ~n238 ;
  assign n240 = x62 ^ x11 ;
  assign n241 = n239 & ~n240 ;
  assign n242 = n236 & ~n241 ;
  assign n243 = x21 ^ x12 ;
  assign n244 = x22 ^ x13 ;
  assign n245 = ~n243 & ~n244 ;
  assign n246 = x23 ^ x14 ;
  assign n247 = n245 & ~n246 ;
  assign n248 = n242 & ~n247 ;
  assign n249 = x24 ^ x12 ;
  assign n250 = x25 ^ x13 ;
  assign n251 = ~n249 & ~n250 ;
  assign n252 = x26 ^ x14 ;
  assign n253 = n251 & ~n252 ;
  assign n254 = n248 & ~n253 ;
  assign n255 = x39 ^ x12 ;
  assign n256 = x40 ^ x13 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = x41 ^ x14 ;
  assign n259 = n257 & ~n258 ;
  assign n260 = n254 & ~n259 ;
  assign n261 = x42 ^ x12 ;
  assign n262 = x43 ^ x13 ;
  assign n263 = ~n261 & ~n262 ;
  assign n264 = x44 ^ x14 ;
  assign n265 = n263 & ~n264 ;
  assign n266 = n260 & ~n265 ;
  assign n267 = x54 ^ x12 ;
  assign n268 = x55 ^ x13 ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = x56 ^ x14 ;
  assign n271 = n269 & ~n270 ;
  assign n272 = n266 & ~n271 ;
  assign n273 = x57 ^ x12 ;
  assign n274 = x58 ^ x13 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = x59 ^ x14 ;
  assign n277 = n275 & ~n276 ;
  assign n278 = n272 & ~n277 ;
  assign n279 = x30 ^ x15 ;
  assign n280 = x31 ^ x16 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = x32 ^ x17 ;
  assign n283 = n281 & ~n282 ;
  assign n284 = n278 & ~n283 ;
  assign n285 = x36 ^ x15 ;
  assign n286 = x37 ^ x16 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = x38 ^ x17 ;
  assign n289 = n287 & ~n288 ;
  assign n290 = n284 & ~n289 ;
  assign n291 = x42 ^ x15 ;
  assign n292 = x43 ^ x16 ;
  assign n293 = ~n291 & ~n292 ;
  assign n294 = x44 ^ x17 ;
  assign n295 = n293 & ~n294 ;
  assign n296 = n290 & ~n295 ;
  assign n297 = x63 ^ x15 ;
  assign n298 = x64 ^ x16 ;
  assign n299 = ~n297 & ~n298 ;
  assign n300 = x65 ^ x17 ;
  assign n301 = n299 & ~n300 ;
  assign n302 = n296 & ~n301 ;
  assign n303 = x30 ^ x18 ;
  assign n304 = x31 ^ x19 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = x32 ^ x20 ;
  assign n307 = n305 & ~n306 ;
  assign n308 = n302 & ~n307 ;
  assign n309 = x33 ^ x18 ;
  assign n310 = x34 ^ x19 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = x35 ^ x20 ;
  assign n313 = n311 & ~n312 ;
  assign n314 = n308 & ~n313 ;
  assign n315 = x39 ^ x18 ;
  assign n316 = x40 ^ x19 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = x41 ^ x20 ;
  assign n319 = n317 & ~n318 ;
  assign n320 = n314 & ~n319 ;
  assign n321 = x63 ^ x18 ;
  assign n322 = x64 ^ x19 ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = x65 ^ x20 ;
  assign n325 = n323 & ~n324 ;
  assign n326 = n320 & ~n325 ;
  assign n327 = x30 ^ x21 ;
  assign n328 = x31 ^ x22 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = x32 ^ x23 ;
  assign n331 = n329 & ~n330 ;
  assign n332 = n326 & ~n331 ;
  assign n333 = x36 ^ x21 ;
  assign n334 = x37 ^ x22 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = x38 ^ x23 ;
  assign n337 = n335 & ~n336 ;
  assign n338 = n332 & ~n337 ;
  assign n339 = x45 ^ x21 ;
  assign n340 = x46 ^ x22 ;
  assign n341 = ~n339 & ~n340 ;
  assign n342 = x47 ^ x23 ;
  assign n343 = n341 & ~n342 ;
  assign n344 = n338 & ~n343 ;
  assign n345 = x63 ^ x21 ;
  assign n346 = x64 ^ x22 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = x65 ^ x23 ;
  assign n349 = n347 & ~n348 ;
  assign n350 = n344 & ~n349 ;
  assign n351 = x30 ^ x24 ;
  assign n352 = x31 ^ x25 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = x32 ^ x26 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = n350 & ~n355 ;
  assign n357 = x33 ^ x24 ;
  assign n358 = x34 ^ x25 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = x35 ^ x26 ;
  assign n361 = n359 & ~n360 ;
  assign n362 = n356 & ~n361 ;
  assign n363 = x45 ^ x24 ;
  assign n364 = x46 ^ x25 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = x47 ^ x26 ;
  assign n367 = n365 & ~n366 ;
  assign n368 = n362 & ~n367 ;
  assign n369 = x63 ^ x24 ;
  assign n370 = x64 ^ x25 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = x65 ^ x26 ;
  assign n373 = n371 & ~n372 ;
  assign n374 = n368 & ~n373 ;
  assign n375 = x30 ^ x27 ;
  assign n376 = x31 ^ x28 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = x32 ^ x29 ;
  assign n379 = n377 & ~n378 ;
  assign n380 = n374 & ~n379 ;
  assign n381 = x39 ^ x27 ;
  assign n382 = x40 ^ x28 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = x41 ^ x29 ;
  assign n385 = n383 & ~n384 ;
  assign n386 = n380 & ~n385 ;
  assign n387 = x42 ^ x27 ;
  assign n388 = x43 ^ x28 ;
  assign n389 = ~n387 & ~n388 ;
  assign n390 = x44 ^ x29 ;
  assign n391 = n389 & ~n390 ;
  assign n392 = n386 & ~n391 ;
  assign n393 = x63 ^ x27 ;
  assign n394 = x64 ^ x28 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = x65 ^ x29 ;
  assign n397 = n395 & ~n396 ;
  assign n398 = n392 & ~n397 ;
  assign n399 = x48 ^ x30 ;
  assign n400 = x49 ^ x31 ;
  assign n401 = ~n399 & ~n400 ;
  assign n402 = x50 ^ x32 ;
  assign n403 = n401 & ~n402 ;
  assign n404 = n398 & ~n403 ;
  assign n405 = x51 ^ x30 ;
  assign n406 = x52 ^ x31 ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = x53 ^ x32 ;
  assign n409 = n407 & ~n408 ;
  assign n410 = n404 & ~n409 ;
  assign n411 = x54 ^ x30 ;
  assign n412 = x55 ^ x31 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = x56 ^ x32 ;
  assign n415 = n413 & ~n414 ;
  assign n416 = n410 & ~n415 ;
  assign n417 = x57 ^ x30 ;
  assign n418 = x58 ^ x31 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = x59 ^ x32 ;
  assign n421 = n419 & ~n420 ;
  assign n422 = n416 & ~n421 ;
  assign n423 = x60 ^ x30 ;
  assign n424 = x61 ^ x31 ;
  assign n425 = ~n423 & ~n424 ;
  assign n426 = x62 ^ x32 ;
  assign n427 = n425 & ~n426 ;
  assign n428 = n422 & ~n427 ;
  assign n429 = x66 ^ x33 ;
  assign n430 = x67 ^ x34 ;
  assign n431 = ~n429 & ~n430 ;
  assign n432 = x68 ^ x35 ;
  assign n433 = n431 & ~n432 ;
  assign n434 = n428 & ~n433 ;
  assign n435 = x66 ^ x36 ;
  assign n436 = x67 ^ x37 ;
  assign n437 = ~n435 & ~n436 ;
  assign n438 = x68 ^ x38 ;
  assign n439 = n437 & ~n438 ;
  assign n440 = n434 & ~n439 ;
  assign n441 = x66 ^ x39 ;
  assign n442 = x67 ^ x40 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = x68 ^ x41 ;
  assign n445 = n443 & ~n444 ;
  assign n446 = n440 & ~n445 ;
  assign n447 = x66 ^ x42 ;
  assign n448 = x67 ^ x43 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = x68 ^ x44 ;
  assign n451 = n449 & ~n450 ;
  assign n452 = n446 & ~n451 ;
  assign n453 = x66 ^ x45 ;
  assign n454 = x67 ^ x46 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = x68 ^ x47 ;
  assign n457 = n455 & ~n456 ;
  assign n458 = n452 & ~n457 ;
  assign n459 = x66 ^ x48 ;
  assign n460 = x67 ^ x49 ;
  assign n461 = ~n459 & ~n460 ;
  assign n462 = x68 ^ x50 ;
  assign n463 = n461 & ~n462 ;
  assign n464 = n458 & ~n463 ;
  assign n465 = x66 ^ x51 ;
  assign n466 = x67 ^ x52 ;
  assign n467 = ~n465 & ~n466 ;
  assign n468 = x68 ^ x53 ;
  assign n469 = n467 & ~n468 ;
  assign n470 = n464 & ~n469 ;
  assign n471 = x66 ^ x54 ;
  assign n472 = x67 ^ x55 ;
  assign n473 = ~n471 & ~n472 ;
  assign n474 = x68 ^ x56 ;
  assign n475 = n473 & ~n474 ;
  assign n476 = n470 & ~n475 ;
  assign n477 = x66 ^ x57 ;
  assign n478 = x67 ^ x58 ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = x68 ^ x59 ;
  assign n481 = n479 & ~n480 ;
  assign n482 = n476 & ~n481 ;
  assign n483 = x66 ^ x60 ;
  assign n484 = x67 ^ x61 ;
  assign n485 = ~n483 & ~n484 ;
  assign n486 = x68 ^ x62 ;
  assign n487 = n485 & ~n486 ;
  assign n488 = n482 & ~n487 ;
  assign n489 = x66 ^ x63 ;
  assign n490 = x67 ^ x64 ;
  assign n491 = ~n489 & ~n490 ;
  assign n492 = x68 ^ x65 ;
  assign n493 = n491 & ~n492 ;
  assign n494 = n488 & ~n493 ;
  assign y0 = n494 ;
endmodule
