module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 ;
  assign n23 = x2 ^ x0 ;
  assign n24 = x3 ^ x1 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = x4 ^ x0 ;
  assign n27 = x5 ^ x1 ;
  assign n28 = ~n26 & ~n27 ;
  assign n29 = ~n25 & ~n28 ;
  assign n30 = x6 ^ x0 ;
  assign n31 = x7 ^ x1 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n29 & ~n32 ;
  assign n34 = x14 ^ x0 ;
  assign n35 = x15 ^ x1 ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = n33 & ~n36 ;
  assign n38 = x6 ^ x2 ;
  assign n39 = x7 ^ x3 ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = n37 & ~n40 ;
  assign n42 = x8 ^ x2 ;
  assign n43 = x9 ^ x3 ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = n41 & ~n44 ;
  assign n46 = x16 ^ x2 ;
  assign n47 = x17 ^ x3 ;
  assign n48 = ~n46 & ~n47 ;
  assign n49 = n45 & ~n48 ;
  assign n50 = x6 ^ x4 ;
  assign n51 = x7 ^ x5 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = n49 & ~n52 ;
  assign n54 = x10 ^ x4 ;
  assign n55 = x11 ^ x5 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = n53 & ~n56 ;
  assign n58 = x12 ^ x4 ;
  assign n59 = x13 ^ x5 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = n57 & ~n60 ;
  assign n62 = x14 ^ x4 ;
  assign n63 = x15 ^ x5 ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = n61 & ~n64 ;
  assign n66 = x18 ^ x4 ;
  assign n67 = x19 ^ x5 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = n65 & ~n68 ;
  assign n70 = x8 ^ x6 ;
  assign n71 = x9 ^ x7 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = n69 & ~n72 ;
  assign n74 = x10 ^ x6 ;
  assign n75 = x11 ^ x7 ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = n73 & ~n76 ;
  assign n78 = x12 ^ x6 ;
  assign n79 = x13 ^ x7 ;
  assign n80 = ~n78 & ~n79 ;
  assign n81 = n77 & ~n80 ;
  assign n82 = x14 ^ x6 ;
  assign n83 = x15 ^ x7 ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = n81 & ~n84 ;
  assign n86 = x12 ^ x8 ;
  assign n87 = x13 ^ x9 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = n85 & ~n88 ;
  assign n90 = x16 ^ x8 ;
  assign n91 = x17 ^ x9 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = n89 & ~n92 ;
  assign n94 = x12 ^ x10 ;
  assign n95 = x13 ^ x11 ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = n93 & ~n96 ;
  assign n98 = x20 ^ x10 ;
  assign n99 = x21 ^ x11 ;
  assign n100 = ~n98 & ~n99 ;
  assign n101 = n97 & ~n100 ;
  assign n102 = x20 ^ x12 ;
  assign n103 = x21 ^ x13 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = n101 & ~n104 ;
  assign n106 = x20 ^ x18 ;
  assign n107 = x21 ^ x19 ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = n105 & ~n108 ;
  assign y0 = n109 ;
endmodule
